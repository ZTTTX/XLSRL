module xls_test(
  input wire clk,
  input wire [511:0] message,
  output wire [255:0] out
);
  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [511:0] p0_message;
  always_ff @ (posedge clk) begin
    p0_message <= message;
  end

  // ===== Pipe stage 1:
  wire [28:0] p1_add_56525_comb;
  wire [30:0] p1_add_56529_comb;
  wire p1_bit_slice_56531_comb;
  wire [31:0] p1_e__66_comb;
  wire [31:0] p1_f__1_comb;
  wire [5:0] p1_S1__67_comb;
  wire [4:0] p1_S1__66_comb;
  wire [13:0] p1_S1__65_comb;
  wire [6:0] p1_S1__64_comb;
  wire [31:0] p1_S1__1_comb;
  wire [31:0] p1_ch__1_comb;
  wire [29:0] p1_add_56559_comb;
  wire [31:0] p1_temp1__336_comb;
  wire [31:0] p1_temp1__337_comb;
  wire [31:0] p1_temp1__338_comb;
  assign p1_add_56525_comb = p0_message[511:483] + 29'h1e6e_fdad;
  assign p1_add_56529_comb = {p1_add_56525_comb, p0_message[482:481]} + 31'h52a7_fa9d;
  assign p1_bit_slice_56531_comb = p0_message[480];
  assign p1_e__66_comb = {p1_add_56529_comb, p1_bit_slice_56531_comb};
  assign p1_f__1_comb = 32'h510e_527f;
  assign p1_S1__67_comb = {p1_add_56529_comb[4:0], p1_bit_slice_56531_comb} ^ p1_add_56529_comb[9:4] ^ p1_add_56529_comb[23:18];
  assign p1_S1__66_comb = p1_add_56529_comb[30:26] ^ {p1_add_56529_comb[3:0], p1_bit_slice_56531_comb} ^ p1_add_56529_comb[17:13];
  assign p1_S1__65_comb = p1_add_56529_comb[25:12] ^ p1_add_56529_comb[30:17] ^ {p1_add_56529_comb[12:0], p1_bit_slice_56531_comb};
  assign p1_S1__64_comb = p1_add_56529_comb[11:5] ^ p1_add_56529_comb[16:10] ^ p1_add_56529_comb[30:24];
  assign p1_S1__1_comb = {p1_S1__67_comb, p1_S1__66_comb, p1_S1__65_comb, p1_S1__64_comb};
  assign p1_ch__1_comb = p1_e__66_comb & p1_f__1_comb ^ ~(p1_e__66_comb | 32'h64fa_9773);
  assign p1_add_56559_comb = p0_message[479:450] + 30'h242e_c78f;
  assign p1_temp1__336_comb = p1_S1__1_comb + p1_ch__1_comb;
  assign p1_temp1__337_comb = {p1_add_56559_comb, p0_message[449:448]};
  assign p1_temp1__338_comb = p1_temp1__336_comb + p1_temp1__337_comb;

  // Registers for pipe stage 1:
  reg [511:0] p1_message;
  reg [28:0] p1_add_56525;
  reg [30:0] p1_add_56529;
  reg p1_bit_slice_56531;
  reg [31:0] p1_e__66;
  reg [31:0] p1_temp1__338;
  always_ff @ (posedge clk) begin
    p1_message <= p0_message;
    p1_add_56525 <= p1_add_56525_comb;
    p1_add_56529 <= p1_add_56529_comb;
    p1_bit_slice_56531 <= p1_bit_slice_56531_comb;
    p1_e__66 <= p1_e__66_comb;
    p1_temp1__338 <= p1_temp1__338_comb;
  end

  // ===== Pipe stage 2:
  wire [30:0] p2_add_56578_comb;
  wire [31:0] p2_e__67_comb;
  wire [5:0] p2_S1__71_comb;
  wire [4:0] p2_S1__70_comb;
  wire [13:0] p2_S1__69_comb;
  wire [6:0] p2_S1__68_comb;
  wire [31:0] p2_S1__2_comb;
  wire [31:0] p2_ch__2_comb;
  wire [31:0] p2_w_im15__1_comb;
  wire [31:0] p2_temp1__331_comb;
  wire [31:0] p2_temp1__332_comb;
  wire [31:0] p2_temp1__333_comb;
  wire [31:0] p2_temp1__334_comb;
  wire [31:0] p2_c__3_comb;
  wire [31:0] p2_e__68_comb;
  wire [2:0] p2_s_0__59_comb;
  wire [3:0] p2_s_0__58_comb;
  wire [10:0] p2_s_0__57_comb;
  wire [13:0] p2_s_0__56_comb;
  wire [31:0] p2_s_0__3_comb;
  wire [31:0] p2_ch__3_comb;
  wire [31:0] p2_concat_56622_comb;
  wire [31:0] p2_value__7_comb;
  assign p2_add_56578_comb = p1_temp1__338[31:1] + 31'h1e37_79b9;
  assign p2_e__67_comb = {p2_add_56578_comb, p1_temp1__338[0]};
  assign p2_S1__71_comb = {p2_add_56578_comb[4:0], p1_temp1__338[0]} ^ p2_add_56578_comb[9:4] ^ p2_add_56578_comb[23:18];
  assign p2_S1__70_comb = p2_add_56578_comb[30:26] ^ {p2_add_56578_comb[3:0], p1_temp1__338[0]} ^ p2_add_56578_comb[17:13];
  assign p2_S1__69_comb = p2_add_56578_comb[25:12] ^ p2_add_56578_comb[30:17] ^ {p2_add_56578_comb[12:0], p1_temp1__338[0]};
  assign p2_S1__68_comb = p2_add_56578_comb[11:5] ^ p2_add_56578_comb[16:10] ^ p2_add_56578_comb[30:24];
  assign p2_S1__2_comb = {p2_S1__71_comb, p2_S1__70_comb, p2_S1__69_comb, p2_S1__68_comb};
  assign p2_ch__2_comb = {p2_add_56578_comb & p1_add_56529, p1_temp1__338[0] & p1_bit_slice_56531} ^ ~(p2_e__67_comb | 32'haef1_ad80);
  assign p2_w_im15__1_comb = p1_message[447:416];
  assign p2_temp1__331_comb = 32'h50c6_645b;
  assign p2_temp1__332_comb = p2_S1__2_comb + p2_ch__2_comb;
  assign p2_temp1__333_comb = p2_w_im15__1_comb + p2_temp1__331_comb;
  assign p2_temp1__334_comb = p2_temp1__332_comb + p2_temp1__333_comb;
  assign p2_c__3_comb = 32'hbb67_ae85;
  assign p2_e__68_comb = p2_temp1__334_comb + p2_c__3_comb;
  assign p2_s_0__59_comb = p1_message[390:388] ^ p1_message[401:399];
  assign p2_s_0__58_comb = p1_message[387:384] ^ p1_message[398:395] ^ p1_message[415:412];
  assign p2_s_0__57_comb = p1_message[415:405] ^ p1_message[394:384] ^ p1_message[411:401];
  assign p2_s_0__56_comb = p1_message[404:391] ^ p1_message[415:402] ^ p1_message[400:387];
  assign p2_s_0__3_comb = {p2_s_0__59_comb, p2_s_0__58_comb, p2_s_0__57_comb, p2_s_0__56_comb};
  assign p2_ch__3_comb = p2_e__68_comb & p2_e__67_comb ^ ~(p2_e__68_comb | {~p1_add_56529, ~p1_bit_slice_56531});
  assign p2_concat_56622_comb = {~p2_add_56578_comb, ~p1_temp1__338[0]};
  assign p2_value__7_comb = p2_w_im15__1_comb + p2_s_0__3_comb;

  // Registers for pipe stage 2:
  reg [511:0] p2_message;
  reg [28:0] p2_add_56525;
  reg [31:0] p2_e__66;
  reg [31:0] p2_temp1__338;
  reg [31:0] p2_e__67;
  reg [31:0] p2_temp1__334;
  reg [31:0] p2_e__68;
  reg [31:0] p2_ch__3;
  reg [31:0] p2_concat_56622;
  reg [31:0] p2_value__7;
  always_ff @ (posedge clk) begin
    p2_message <= p1_message;
    p2_add_56525 <= p1_add_56525;
    p2_e__66 <= p1_e__66;
    p2_temp1__338 <= p1_temp1__338;
    p2_e__67 <= p2_e__67_comb;
    p2_temp1__334 <= p2_temp1__334_comb;
    p2_e__68 <= p2_e__68_comb;
    p2_ch__3 <= p2_ch__3_comb;
    p2_concat_56622 <= p2_concat_56622_comb;
    p2_value__7 <= p2_value__7_comb;
  end

  // ===== Pipe stage 3:
  wire [5:0] p3_S1__75_comb;
  wire [4:0] p3_S1__74_comb;
  wire [13:0] p3_S1__73_comb;
  wire [6:0] p3_S1__72_comb;
  wire [31:0] p3_S1__3_comb;
  wire [29:0] p3_add_56679_comb;
  wire [31:0] p3_temp1__328_comb;
  wire [31:0] p3_temp1__329_comb;
  wire [31:0] p3_temp1__323_comb;
  wire [31:0] p3_temp2_comb;
  wire [31:0] p3_temp1__330_comb;
  wire [31:0] p3_b__3_comb;
  wire [31:0] p3_a__1_comb;
  wire [31:0] p3_e__69_comb;
  wire [31:0] p3_b__67_comb;
  wire [31:0] p3_c__67_comb;
  wire [1:0] p3_S0__67_comb;
  wire [10:0] p3_S0__66_comb;
  wire [8:0] p3_S0__65_comb;
  wire [9:0] p3_S0__64_comb;
  wire [31:0] p3_and_56729_comb;
  wire [5:0] p3_S1__79_comb;
  wire [4:0] p3_S1__78_comb;
  wire [13:0] p3_S1__77_comb;
  wire [6:0] p3_S1__76_comb;
  wire [31:0] p3_S0__1_comb;
  wire [31:0] p3_maj__1_comb;
  wire [31:0] p3_S1__4_comb;
  wire [31:0] p3_temp2__1_comb;
  wire [31:0] p3_temp1__17_comb;
  wire [31:0] p3_ch__4_comb;
  wire [31:0] p3_a__2_comb;
  assign p3_S1__75_comb = p2_e__68[5:0] ^ p2_e__68[10:5] ^ p2_e__68[24:19];
  assign p3_S1__74_comb = p2_e__68[31:27] ^ p2_e__68[4:0] ^ p2_e__68[18:14];
  assign p3_S1__73_comb = p2_e__68[26:13] ^ p2_e__68[31:18] ^ p2_e__68[13:0];
  assign p3_S1__72_comb = p2_e__68[12:6] ^ p2_e__68[17:11] ^ p2_e__68[31:25];
  assign p3_S1__3_comb = {p3_S1__75_comb, p3_S1__74_comb, p3_S1__73_comb, p3_S1__72_comb};
  assign p3_add_56679_comb = p2_message[415:386] + 30'h0eb1_0b89;
  assign p3_temp1__328_comb = p3_S1__3_comb + p2_ch__3;
  assign p3_temp1__329_comb = {p3_add_56679_comb, p2_message[385:384]};
  assign p3_temp1__323_comb = {p2_add_56525, p2_message[482:480]};
  assign p3_temp2_comb = 32'h0890_9ae5;
  assign p3_temp1__330_comb = p3_temp1__328_comb + p3_temp1__329_comb;
  assign p3_b__3_comb = 32'h6a09_e667;
  assign p3_a__1_comb = p3_temp1__323_comb + p3_temp2_comb;
  assign p3_e__69_comb = p3_temp1__330_comb + p3_b__3_comb;
  assign p3_b__67_comb = 32'h6a09_e667;
  assign p3_c__67_comb = 32'hbb67_ae85;
  assign p3_S0__67_comb = p3_a__1_comb[1:0] ^ p3_a__1_comb[12:11] ^ p3_a__1_comb[21:20];
  assign p3_S0__66_comb = p3_a__1_comb[31:21] ^ p3_a__1_comb[10:0] ^ p3_a__1_comb[19:9];
  assign p3_S0__65_comb = p3_a__1_comb[20:12] ^ p3_a__1_comb[31:23] ^ p3_a__1_comb[8:0];
  assign p3_S0__64_comb = p3_a__1_comb[11:2] ^ p3_a__1_comb[22:13] ^ p3_a__1_comb[31:22];
  assign p3_and_56729_comb = p3_a__1_comb & p3_b__67_comb;
  assign p3_S1__79_comb = p3_e__69_comb[5:0] ^ p3_e__69_comb[10:5] ^ p3_e__69_comb[24:19];
  assign p3_S1__78_comb = p3_e__69_comb[31:27] ^ p3_e__69_comb[4:0] ^ p3_e__69_comb[18:14];
  assign p3_S1__77_comb = p3_e__69_comb[26:13] ^ p3_e__69_comb[31:18] ^ p3_e__69_comb[13:0];
  assign p3_S1__76_comb = p3_e__69_comb[12:6] ^ p3_e__69_comb[17:11] ^ p3_e__69_comb[31:25];
  assign p3_S0__1_comb = {p3_S0__67_comb, p3_S0__66_comb, p3_S0__65_comb, p3_S0__64_comb};
  assign p3_maj__1_comb = p3_and_56729_comb ^ p3_a__1_comb & p3_c__67_comb ^ 32'h2a01_a605;
  assign p3_S1__4_comb = {p3_S1__79_comb, p3_S1__78_comb, p3_S1__77_comb, p3_S1__76_comb};
  assign p3_temp2__1_comb = p3_S0__1_comb + p3_maj__1_comb;
  assign p3_temp1__17_comb = p2_e__66 + p3_S1__4_comb;
  assign p3_ch__4_comb = p3_e__69_comb & p2_e__68 ^ ~(p3_e__69_comb | p2_concat_56622);
  assign p3_a__2_comb = p2_temp1__338 + p3_temp2__1_comb;

  // Registers for pipe stage 3:
  reg [511:0] p3_message;
  reg [31:0] p3_e__67;
  reg [31:0] p3_temp1__334;
  reg [31:0] p3_e__68;
  reg [31:0] p3_temp1__330;
  reg [31:0] p3_e__69;
  reg [31:0] p3_temp1__17;
  reg [31:0] p3_ch__4;
  reg [31:0] p3_a__1;
  reg [31:0] p3_and_56729;
  reg [31:0] p3_a__2;
  reg [31:0] p3_value__7;
  always_ff @ (posedge clk) begin
    p3_message <= p2_message;
    p3_e__67 <= p2_e__67;
    p3_temp1__334 <= p2_temp1__334;
    p3_e__68 <= p2_e__68;
    p3_temp1__330 <= p3_temp1__330_comb;
    p3_e__69 <= p3_e__69_comb;
    p3_temp1__17 <= p3_temp1__17_comb;
    p3_ch__4 <= p3_ch__4_comb;
    p3_a__1 <= p3_a__1_comb;
    p3_and_56729 <= p3_and_56729_comb;
    p3_a__2 <= p3_a__2_comb;
    p3_value__7 <= p2_value__7;
  end

  // ===== Pipe stage 4:
  wire [31:0] p4_b__2_comb;
  wire [1:0] p4_S0__71_comb;
  wire [10:0] p4_S0__70_comb;
  wire [8:0] p4_S0__69_comb;
  wire [9:0] p4_S0__68_comb;
  wire [31:0] p4_and_56801_comb;
  wire [31:0] p4_w_im15__3_comb;
  wire [31:0] p4_S0__2_comb;
  wire [31:0] p4_maj__2_comb;
  wire [31:0] p4_temp1__18_comb;
  wire [31:0] p4_temp1__262_comb;
  wire [31:0] p4_temp2__2_comb;
  wire [31:0] p4_temp1__20_comb;
  wire [31:0] p4_a__3_comb;
  wire [31:0] p4_e__5_comb;
  wire [1:0] p4_S0__75_comb;
  wire [10:0] p4_S0__74_comb;
  wire [8:0] p4_S0__73_comb;
  wire [9:0] p4_S0__72_comb;
  wire [31:0] p4_and_56823_comb;
  wire [5:0] p4_S1__83_comb;
  wire [4:0] p4_S1__82_comb;
  wire [13:0] p4_S1__81_comb;
  wire [6:0] p4_S1__80_comb;
  wire [31:0] p4_S0__3_comb;
  wire [31:0] p4_maj__3_comb;
  wire [2:0] p4_s_0__67_comb;
  wire [3:0] p4_s_0__66_comb;
  wire [10:0] p4_s_0__65_comb;
  wire [13:0] p4_s_0__64_comb;
  wire [31:0] p4_S1__5_comb;
  wire [31:0] p4_temp2__3_comb;
  wire [31:0] p4_s_0__5_comb;
  wire [31:0] p4_temp1__21_comb;
  wire [31:0] p4_a__4_comb;
  wire [31:0] p4_value__13_comb;
  assign p4_b__2_comb = 32'h6a09_e667;
  assign p4_S0__71_comb = p3_a__2[1:0] ^ p3_a__2[12:11] ^ p3_a__2[21:20];
  assign p4_S0__70_comb = p3_a__2[31:21] ^ p3_a__2[10:0] ^ p3_a__2[19:9];
  assign p4_S0__69_comb = p3_a__2[20:12] ^ p3_a__2[31:23] ^ p3_a__2[8:0];
  assign p4_S0__68_comb = p3_a__2[11:2] ^ p3_a__2[22:13] ^ p3_a__2[31:22];
  assign p4_and_56801_comb = p3_a__2 & p3_a__1;
  assign p4_w_im15__3_comb = p3_message[383:352];
  assign p4_S0__2_comb = {p4_S0__71_comb, p4_S0__70_comb, p4_S0__69_comb, p4_S0__68_comb};
  assign p4_maj__2_comb = p4_and_56801_comb ^ p3_a__2 & p4_b__2_comb ^ p3_and_56729;
  assign p4_temp1__18_comb = p3_temp1__17 + p3_ch__4;
  assign p4_temp1__262_comb = p4_w_im15__3_comb + 32'h3956_c25b;
  assign p4_temp2__2_comb = p4_S0__2_comb + p4_maj__2_comb;
  assign p4_temp1__20_comb = p4_temp1__18_comb + p4_temp1__262_comb;
  assign p4_a__3_comb = p3_temp1__334 + p4_temp2__2_comb;
  assign p4_e__5_comb = p3_a__1 + p4_temp1__20_comb;
  assign p4_S0__75_comb = p4_a__3_comb[1:0] ^ p4_a__3_comb[12:11] ^ p4_a__3_comb[21:20];
  assign p4_S0__74_comb = p4_a__3_comb[31:21] ^ p4_a__3_comb[10:0] ^ p4_a__3_comb[19:9];
  assign p4_S0__73_comb = p4_a__3_comb[20:12] ^ p4_a__3_comb[31:23] ^ p4_a__3_comb[8:0];
  assign p4_S0__72_comb = p4_a__3_comb[11:2] ^ p4_a__3_comb[22:13] ^ p4_a__3_comb[31:22];
  assign p4_and_56823_comb = p4_a__3_comb & p3_a__2;
  assign p4_S1__83_comb = p4_e__5_comb[5:0] ^ p4_e__5_comb[10:5] ^ p4_e__5_comb[24:19];
  assign p4_S1__82_comb = p4_e__5_comb[31:27] ^ p4_e__5_comb[4:0] ^ p4_e__5_comb[18:14];
  assign p4_S1__81_comb = p4_e__5_comb[26:13] ^ p4_e__5_comb[31:18] ^ p4_e__5_comb[13:0];
  assign p4_S1__80_comb = p4_e__5_comb[12:6] ^ p4_e__5_comb[17:11] ^ p4_e__5_comb[31:25];
  assign p4_S0__3_comb = {p4_S0__75_comb, p4_S0__74_comb, p4_S0__73_comb, p4_S0__72_comb};
  assign p4_maj__3_comb = p4_and_56823_comb ^ p4_a__3_comb & p3_a__1 ^ p4_and_56801_comb;
  assign p4_s_0__67_comb = p3_message[326:324] ^ p3_message[337:335];
  assign p4_s_0__66_comb = p3_message[323:320] ^ p3_message[334:331] ^ p3_message[351:348];
  assign p4_s_0__65_comb = p3_message[351:341] ^ p3_message[330:320] ^ p3_message[347:337];
  assign p4_s_0__64_comb = p3_message[340:327] ^ p3_message[351:338] ^ p3_message[336:323];
  assign p4_S1__5_comb = {p4_S1__83_comb, p4_S1__82_comb, p4_S1__81_comb, p4_S1__80_comb};
  assign p4_temp2__3_comb = p4_S0__3_comb + p4_maj__3_comb;
  assign p4_s_0__5_comb = {p4_s_0__67_comb, p4_s_0__66_comb, p4_s_0__65_comb, p4_s_0__64_comb};
  assign p4_temp1__21_comb = p3_e__67 + p4_S1__5_comb;
  assign p4_a__4_comb = p3_temp1__330 + p4_temp2__3_comb;
  assign p4_value__13_comb = p4_w_im15__3_comb + p4_s_0__5_comb;

  // Registers for pipe stage 4:
  reg [511:0] p4_message;
  reg [31:0] p4_e__68;
  reg [31:0] p4_e__69;
  reg [31:0] p4_temp1__20;
  reg [31:0] p4_e__5;
  reg [31:0] p4_temp1__21;
  reg [31:0] p4_a__2;
  reg [31:0] p4_a__3;
  reg [31:0] p4_and_56823;
  reg [31:0] p4_a__4;
  reg [31:0] p4_value__7;
  reg [31:0] p4_value__13;
  always_ff @ (posedge clk) begin
    p4_message <= p3_message;
    p4_e__68 <= p3_e__68;
    p4_e__69 <= p3_e__69;
    p4_temp1__20 <= p4_temp1__20_comb;
    p4_e__5 <= p4_e__5_comb;
    p4_temp1__21 <= p4_temp1__21_comb;
    p4_a__2 <= p3_a__2;
    p4_a__3 <= p4_a__3_comb;
    p4_and_56823 <= p4_and_56823_comb;
    p4_a__4 <= p4_a__4_comb;
    p4_value__7 <= p3_value__7;
    p4_value__13 <= p4_value__13_comb;
  end

  // ===== Pipe stage 5:
  wire [1:0] p5_S0__79_comb;
  wire [10:0] p5_S0__78_comb;
  wire [8:0] p5_S0__77_comb;
  wire [9:0] p5_S0__76_comb;
  wire [31:0] p5_and_56924_comb;
  wire [31:0] p5_ch__5_comb;
  wire [31:0] p5_w_im15__4_comb;
  wire [31:0] p5_S0__4_comb;
  wire [31:0] p5_maj__4_comb;
  wire [31:0] p5_temp1__22_comb;
  wire [31:0] p5_temp1__263_comb;
  wire [31:0] p5_temp2__4_comb;
  wire [31:0] p5_temp1__24_comb;
  wire [31:0] p5_a__5_comb;
  wire [31:0] p5_e__6_comb;
  wire [1:0] p5_S0__83_comb;
  wire [10:0] p5_S0__82_comb;
  wire [8:0] p5_S0__81_comb;
  wire [9:0] p5_S0__80_comb;
  wire [31:0] p5_and_56946_comb;
  wire [5:0] p5_S1__87_comb;
  wire [4:0] p5_S1__86_comb;
  wire [13:0] p5_S1__85_comb;
  wire [6:0] p5_S1__84_comb;
  wire [29:0] p5_add_56901_comb;
  wire [31:0] p5_S0__5_comb;
  wire [31:0] p5_maj__5_comb;
  wire [2:0] p5_s_0__71_comb;
  wire [3:0] p5_s_0__70_comb;
  wire [10:0] p5_s_0__69_comb;
  wire [13:0] p5_s_0__68_comb;
  wire [31:0] p5_S1__6_comb;
  wire [31:0] p5_ch__6_comb;
  wire [31:0] p5_temp1__264_comb;
  wire [31:0] p5_temp2__5_comb;
  wire [31:0] p5_s_0__6_comb;
  wire [31:0] p5_temp1__437_comb;
  wire [31:0] p5_temp1__438_comb;
  wire [31:0] p5_a__6_comb;
  wire [31:0] p5_value__16_comb;
  assign p5_S0__79_comb = p4_a__4[1:0] ^ p4_a__4[12:11] ^ p4_a__4[21:20];
  assign p5_S0__78_comb = p4_a__4[31:21] ^ p4_a__4[10:0] ^ p4_a__4[19:9];
  assign p5_S0__77_comb = p4_a__4[20:12] ^ p4_a__4[31:23] ^ p4_a__4[8:0];
  assign p5_S0__76_comb = p4_a__4[11:2] ^ p4_a__4[22:13] ^ p4_a__4[31:22];
  assign p5_and_56924_comb = p4_a__4 & p4_a__3;
  assign p5_ch__5_comb = p4_e__5 & p4_e__69 ^ ~(p4_e__5 | ~p4_e__68);
  assign p5_w_im15__4_comb = p4_message[351:320];
  assign p5_S0__4_comb = {p5_S0__79_comb, p5_S0__78_comb, p5_S0__77_comb, p5_S0__76_comb};
  assign p5_maj__4_comb = p5_and_56924_comb ^ p4_a__4 & p4_a__2 ^ p4_and_56823;
  assign p5_temp1__22_comb = p4_temp1__21 + p5_ch__5_comb;
  assign p5_temp1__263_comb = p5_w_im15__4_comb + 32'h59f1_11f1;
  assign p5_temp2__4_comb = p5_S0__4_comb + p5_maj__4_comb;
  assign p5_temp1__24_comb = p5_temp1__22_comb + p5_temp1__263_comb;
  assign p5_a__5_comb = p4_temp1__20 + p5_temp2__4_comb;
  assign p5_e__6_comb = p4_a__2 + p5_temp1__24_comb;
  assign p5_S0__83_comb = p5_a__5_comb[1:0] ^ p5_a__5_comb[12:11] ^ p5_a__5_comb[21:20];
  assign p5_S0__82_comb = p5_a__5_comb[31:21] ^ p5_a__5_comb[10:0] ^ p5_a__5_comb[19:9];
  assign p5_S0__81_comb = p5_a__5_comb[20:12] ^ p5_a__5_comb[31:23] ^ p5_a__5_comb[8:0];
  assign p5_S0__80_comb = p5_a__5_comb[11:2] ^ p5_a__5_comb[22:13] ^ p5_a__5_comb[31:22];
  assign p5_and_56946_comb = p5_a__5_comb & p4_a__4;
  assign p5_S1__87_comb = p5_e__6_comb[5:0] ^ p5_e__6_comb[10:5] ^ p5_e__6_comb[24:19];
  assign p5_S1__86_comb = p5_e__6_comb[31:27] ^ p5_e__6_comb[4:0] ^ p5_e__6_comb[18:14];
  assign p5_S1__85_comb = p5_e__6_comb[26:13] ^ p5_e__6_comb[31:18] ^ p5_e__6_comb[13:0];
  assign p5_S1__84_comb = p5_e__6_comb[12:6] ^ p5_e__6_comb[17:11] ^ p5_e__6_comb[31:25];
  assign p5_add_56901_comb = p4_message[319:290] + 30'h248f_e0a9;
  assign p5_S0__5_comb = {p5_S0__83_comb, p5_S0__82_comb, p5_S0__81_comb, p5_S0__80_comb};
  assign p5_maj__5_comb = p5_and_56946_comb ^ p5_a__5_comb & p4_a__3 ^ p5_and_56924_comb;
  assign p5_s_0__71_comb = p4_message[294:292] ^ p4_message[305:303];
  assign p5_s_0__70_comb = p4_message[291:288] ^ p4_message[302:299] ^ p4_message[319:316];
  assign p5_s_0__69_comb = p4_message[319:309] ^ p4_message[298:288] ^ p4_message[315:305];
  assign p5_s_0__68_comb = p4_message[308:295] ^ p4_message[319:306] ^ p4_message[304:291];
  assign p5_S1__6_comb = {p5_S1__87_comb, p5_S1__86_comb, p5_S1__85_comb, p5_S1__84_comb};
  assign p5_ch__6_comb = p5_e__6_comb & p4_e__5 ^ ~(p5_e__6_comb | ~p4_e__69);
  assign p5_temp1__264_comb = {p5_add_56901_comb, p4_message[289:288]};
  assign p5_temp2__5_comb = p5_S0__5_comb + p5_maj__5_comb;
  assign p5_s_0__6_comb = {p5_s_0__71_comb, p5_s_0__70_comb, p5_s_0__69_comb, p5_s_0__68_comb};
  assign p5_temp1__437_comb = p4_e__68 + p5_S1__6_comb;
  assign p5_temp1__438_comb = p5_ch__6_comb + p5_temp1__264_comb;
  assign p5_a__6_comb = p5_temp1__24_comb + p5_temp2__5_comb;
  assign p5_value__16_comb = p5_w_im15__4_comb + p5_s_0__6_comb;

  // Registers for pipe stage 5:
  reg [511:0] p5_message;
  reg [31:0] p5_e__69;
  reg [31:0] p5_e__5;
  reg [31:0] p5_e__6;
  reg [31:0] p5_temp1__437;
  reg [31:0] p5_temp1__438;
  reg [31:0] p5_a__3;
  reg [31:0] p5_a__4;
  reg [31:0] p5_a__5;
  reg [31:0] p5_and_56946;
  reg [31:0] p5_a__6;
  reg [31:0] p5_value__7;
  reg [31:0] p5_value__13;
  reg [31:0] p5_value__16;
  always_ff @ (posedge clk) begin
    p5_message <= p4_message;
    p5_e__69 <= p4_e__69;
    p5_e__5 <= p4_e__5;
    p5_e__6 <= p5_e__6_comb;
    p5_temp1__437 <= p5_temp1__437_comb;
    p5_temp1__438 <= p5_temp1__438_comb;
    p5_a__3 <= p4_a__3;
    p5_a__4 <= p4_a__4;
    p5_a__5 <= p5_a__5_comb;
    p5_and_56946 <= p5_and_56946_comb;
    p5_a__6 <= p5_a__6_comb;
    p5_value__7 <= p4_value__7;
    p5_value__13 <= p4_value__13;
    p5_value__16 <= p5_value__16_comb;
  end

  // ===== Pipe stage 6:
  wire [31:0] p6_temp1__439_comb;
  wire [31:0] p6_e__7_comb;
  wire [5:0] p6_S1__91_comb;
  wire [4:0] p6_S1__90_comb;
  wire [13:0] p6_S1__89_comb;
  wire [6:0] p6_S1__88_comb;
  wire [1:0] p6_S0__87_comb;
  wire [10:0] p6_S0__86_comb;
  wire [8:0] p6_S0__85_comb;
  wire [9:0] p6_S0__84_comb;
  wire [31:0] p6_and_57041_comb;
  wire [31:0] p6_S1__7_comb;
  wire [31:0] p6_S0__6_comb;
  wire [31:0] p6_maj__6_comb;
  wire [2:0] p6_s_0__79_comb;
  wire [3:0] p6_s_0__78_comb;
  wire [10:0] p6_s_0__77_comb;
  wire [13:0] p6_s_0__76_comb;
  wire [31:0] p6_temp1__29_comb;
  wire [31:0] p6_ch__7_comb;
  wire [31:0] p6_w_im15__6_comb;
  wire [31:0] p6_temp2__6_comb;
  wire [31:0] p6_s_0__8_comb;
  wire [31:0] p6_temp1__30_comb;
  wire [31:0] p6_temp1__265_comb;
  wire [31:0] p6_a__7_comb;
  wire [31:0] p6_value__22_comb;
  assign p6_temp1__439_comb = p5_temp1__437 + p5_temp1__438;
  assign p6_e__7_comb = p5_a__3 + p6_temp1__439_comb;
  assign p6_S1__91_comb = p6_e__7_comb[5:0] ^ p6_e__7_comb[10:5] ^ p6_e__7_comb[24:19];
  assign p6_S1__90_comb = p6_e__7_comb[31:27] ^ p6_e__7_comb[4:0] ^ p6_e__7_comb[18:14];
  assign p6_S1__89_comb = p6_e__7_comb[26:13] ^ p6_e__7_comb[31:18] ^ p6_e__7_comb[13:0];
  assign p6_S1__88_comb = p6_e__7_comb[12:6] ^ p6_e__7_comb[17:11] ^ p6_e__7_comb[31:25];
  assign p6_S0__87_comb = p5_a__6[1:0] ^ p5_a__6[12:11] ^ p5_a__6[21:20];
  assign p6_S0__86_comb = p5_a__6[31:21] ^ p5_a__6[10:0] ^ p5_a__6[19:9];
  assign p6_S0__85_comb = p5_a__6[20:12] ^ p5_a__6[31:23] ^ p5_a__6[8:0];
  assign p6_S0__84_comb = p5_a__6[11:2] ^ p5_a__6[22:13] ^ p5_a__6[31:22];
  assign p6_and_57041_comb = p5_a__6 & p5_a__5;
  assign p6_S1__7_comb = {p6_S1__91_comb, p6_S1__90_comb, p6_S1__89_comb, p6_S1__88_comb};
  assign p6_S0__6_comb = {p6_S0__87_comb, p6_S0__86_comb, p6_S0__85_comb, p6_S0__84_comb};
  assign p6_maj__6_comb = p6_and_57041_comb ^ p5_a__6 & p5_a__4 ^ p5_and_56946;
  assign p6_s_0__79_comb = p5_message[230:228] ^ p5_message[241:239];
  assign p6_s_0__78_comb = p5_message[227:224] ^ p5_message[238:235] ^ p5_message[255:252];
  assign p6_s_0__77_comb = p5_message[255:245] ^ p5_message[234:224] ^ p5_message[251:241];
  assign p6_s_0__76_comb = p5_message[244:231] ^ p5_message[255:242] ^ p5_message[240:227];
  assign p6_temp1__29_comb = p5_e__69 + p6_S1__7_comb;
  assign p6_ch__7_comb = p6_e__7_comb & p5_e__6 ^ ~(p6_e__7_comb | ~p5_e__5);
  assign p6_w_im15__6_comb = p5_message[287:256];
  assign p6_temp2__6_comb = p6_S0__6_comb + p6_maj__6_comb;
  assign p6_s_0__8_comb = {p6_s_0__79_comb, p6_s_0__78_comb, p6_s_0__77_comb, p6_s_0__76_comb};
  assign p6_temp1__30_comb = p6_temp1__29_comb + p6_ch__7_comb;
  assign p6_temp1__265_comb = p6_w_im15__6_comb + 32'hab1c_5ed5;
  assign p6_a__7_comb = p6_temp1__439_comb + p6_temp2__6_comb;
  assign p6_value__22_comb = p6_w_im15__6_comb + p6_s_0__8_comb;

  // Registers for pipe stage 6:
  reg [511:0] p6_message;
  reg [31:0] p6_e__5;
  reg [31:0] p6_e__6;
  reg [31:0] p6_e__7;
  reg [31:0] p6_temp1__30;
  reg [31:0] p6_temp1__265;
  reg [31:0] p6_a__4;
  reg [31:0] p6_a__5;
  reg [31:0] p6_a__6;
  reg [31:0] p6_and_57041;
  reg [31:0] p6_a__7;
  reg [31:0] p6_value__7;
  reg [31:0] p6_value__13;
  reg [31:0] p6_value__16;
  reg [31:0] p6_value__22;
  always_ff @ (posedge clk) begin
    p6_message <= p5_message;
    p6_e__5 <= p5_e__5;
    p6_e__6 <= p5_e__6;
    p6_e__7 <= p6_e__7_comb;
    p6_temp1__30 <= p6_temp1__30_comb;
    p6_temp1__265 <= p6_temp1__265_comb;
    p6_a__4 <= p5_a__4;
    p6_a__5 <= p5_a__5;
    p6_a__6 <= p5_a__6;
    p6_and_57041 <= p6_and_57041_comb;
    p6_a__7 <= p6_a__7_comb;
    p6_value__7 <= p5_value__7;
    p6_value__13 <= p5_value__13;
    p6_value__16 <= p5_value__16;
    p6_value__22 <= p6_value__22_comb;
  end

  // ===== Pipe stage 7:
  wire [31:0] p7_temp1__32_comb;
  wire [31:0] p7_e__8_comb;
  wire [5:0] p7_S1__95_comb;
  wire [4:0] p7_S1__94_comb;
  wire [13:0] p7_S1__93_comb;
  wire [6:0] p7_S1__92_comb;
  wire [28:0] p7_add_57117_comb;
  wire [1:0] p7_S0__91_comb;
  wire [10:0] p7_S0__90_comb;
  wire [8:0] p7_S0__89_comb;
  wire [9:0] p7_S0__88_comb;
  wire [31:0] p7_and_57141_comb;
  wire [31:0] p7_S1__8_comb;
  wire [31:0] p7_ch__8_comb;
  wire [31:0] p7_temp1__266_comb;
  wire [31:0] p7_S0__7_comb;
  wire [31:0] p7_maj__7_comb;
  wire [31:0] p7_temp1__434_comb;
  wire [31:0] p7_temp1__435_comb;
  wire [31:0] p7_temp2__7_comb;
  wire [31:0] p7_temp1__436_comb;
  wire [31:0] p7_a__8_comb;
  assign p7_temp1__32_comb = p6_temp1__30 + p6_temp1__265;
  assign p7_e__8_comb = p6_a__4 + p7_temp1__32_comb;
  assign p7_S1__95_comb = p7_e__8_comb[5:0] ^ p7_e__8_comb[10:5] ^ p7_e__8_comb[24:19];
  assign p7_S1__94_comb = p7_e__8_comb[31:27] ^ p7_e__8_comb[4:0] ^ p7_e__8_comb[18:14];
  assign p7_S1__93_comb = p7_e__8_comb[26:13] ^ p7_e__8_comb[31:18] ^ p7_e__8_comb[13:0];
  assign p7_S1__92_comb = p7_e__8_comb[12:6] ^ p7_e__8_comb[17:11] ^ p7_e__8_comb[31:25];
  assign p7_add_57117_comb = p6_message[255:227] + 29'h1b00_f553;
  assign p7_S0__91_comb = p6_a__7[1:0] ^ p6_a__7[12:11] ^ p6_a__7[21:20];
  assign p7_S0__90_comb = p6_a__7[31:21] ^ p6_a__7[10:0] ^ p6_a__7[19:9];
  assign p7_S0__89_comb = p6_a__7[20:12] ^ p6_a__7[31:23] ^ p6_a__7[8:0];
  assign p7_S0__88_comb = p6_a__7[11:2] ^ p6_a__7[22:13] ^ p6_a__7[31:22];
  assign p7_and_57141_comb = p6_a__7 & p6_a__6;
  assign p7_S1__8_comb = {p7_S1__95_comb, p7_S1__94_comb, p7_S1__93_comb, p7_S1__92_comb};
  assign p7_ch__8_comb = p7_e__8_comb & p6_e__7 ^ ~(p7_e__8_comb | ~p6_e__6);
  assign p7_temp1__266_comb = {p7_add_57117_comb, p6_message[226:224]};
  assign p7_S0__7_comb = {p7_S0__91_comb, p7_S0__90_comb, p7_S0__89_comb, p7_S0__88_comb};
  assign p7_maj__7_comb = p7_and_57141_comb ^ p6_a__7 & p6_a__5 ^ p6_and_57041;
  assign p7_temp1__434_comb = p6_e__5 + p7_S1__8_comb;
  assign p7_temp1__435_comb = p7_ch__8_comb + p7_temp1__266_comb;
  assign p7_temp2__7_comb = p7_S0__7_comb + p7_maj__7_comb;
  assign p7_temp1__436_comb = p7_temp1__434_comb + p7_temp1__435_comb;
  assign p7_a__8_comb = p7_temp1__32_comb + p7_temp2__7_comb;

  // Registers for pipe stage 7:
  reg [511:0] p7_message;
  reg [31:0] p7_e__6;
  reg [31:0] p7_e__7;
  reg [31:0] p7_e__8;
  reg [31:0] p7_a__5;
  reg [31:0] p7_temp1__436;
  reg [31:0] p7_a__6;
  reg [31:0] p7_a__7;
  reg [31:0] p7_and_57141;
  reg [31:0] p7_a__8;
  reg [31:0] p7_value__7;
  reg [31:0] p7_value__13;
  reg [31:0] p7_value__16;
  reg [31:0] p7_value__22;
  always_ff @ (posedge clk) begin
    p7_message <= p6_message;
    p7_e__6 <= p6_e__6;
    p7_e__7 <= p6_e__7;
    p7_e__8 <= p7_e__8_comb;
    p7_a__5 <= p6_a__5;
    p7_temp1__436 <= p7_temp1__436_comb;
    p7_a__6 <= p6_a__6;
    p7_a__7 <= p6_a__7;
    p7_and_57141 <= p7_and_57141_comb;
    p7_a__8 <= p7_a__8_comb;
    p7_value__7 <= p6_value__7;
    p7_value__13 <= p6_value__13;
    p7_value__16 <= p6_value__16;
    p7_value__22 <= p6_value__22;
  end

  // ===== Pipe stage 8:
  wire [31:0] p8_e__9_comb;
  wire [5:0] p8_S1__99_comb;
  wire [4:0] p8_S1__98_comb;
  wire [13:0] p8_S1__97_comb;
  wire [6:0] p8_S1__96_comb;
  wire [31:0] p8_S1__9_comb;
  wire [1:0] p8_S0__95_comb;
  wire [10:0] p8_S0__94_comb;
  wire [8:0] p8_S0__93_comb;
  wire [9:0] p8_S0__92_comb;
  wire [31:0] p8_and_57219_comb;
  wire [2:0] p8_s_0__51_comb;
  wire [3:0] p8_s_0__50_comb;
  wire [10:0] p8_s_0__49_comb;
  wire [13:0] p8_s_0__48_comb;
  wire [9:0] p8_s_1__51_comb;
  wire [6:0] p8_s_1__50_comb;
  wire [1:0] p8_s_1__49_comb;
  wire [12:0] p8_s_1__48_comb;
  wire [31:0] p8_temp1__37_comb;
  wire [31:0] p8_ch__9_comb;
  wire [31:0] p8_w_im15__8_comb;
  wire [31:0] p8_S0__8_comb;
  wire [31:0] p8_maj__8_comb;
  wire [31:0] p8_s_0__1_comb;
  wire [31:0] p8_s_1__1_comb;
  wire [2:0] p8_s_0__87_comb;
  wire [3:0] p8_s_0__86_comb;
  wire [10:0] p8_s_0__85_comb;
  wire [13:0] p8_s_0__84_comb;
  wire [31:0] p8_temp1__38_comb;
  wire [31:0] p8_temp1__267_comb;
  wire [31:0] p8_temp2__8_comb;
  wire [31:0] p8_value__1_comb;
  wire [31:0] p8_value__2_comb;
  wire [31:0] p8_s_0__10_comb;
  wire [31:0] p8_temp1__40_comb;
  wire [31:0] p8_a__9_comb;
  wire [31:0] p8_value__3_comb;
  wire [31:0] p8_value__28_comb;
  assign p8_e__9_comb = p7_a__5 + p7_temp1__436;
  assign p8_S1__99_comb = p8_e__9_comb[5:0] ^ p8_e__9_comb[10:5] ^ p8_e__9_comb[24:19];
  assign p8_S1__98_comb = p8_e__9_comb[31:27] ^ p8_e__9_comb[4:0] ^ p8_e__9_comb[18:14];
  assign p8_S1__97_comb = p8_e__9_comb[26:13] ^ p8_e__9_comb[31:18] ^ p8_e__9_comb[13:0];
  assign p8_S1__96_comb = p8_e__9_comb[12:6] ^ p8_e__9_comb[17:11] ^ p8_e__9_comb[31:25];
  assign p8_S1__9_comb = {p8_S1__99_comb, p8_S1__98_comb, p8_S1__97_comb, p8_S1__96_comb};
  assign p8_S0__95_comb = p7_a__8[1:0] ^ p7_a__8[12:11] ^ p7_a__8[21:20];
  assign p8_S0__94_comb = p7_a__8[31:21] ^ p7_a__8[10:0] ^ p7_a__8[19:9];
  assign p8_S0__93_comb = p7_a__8[20:12] ^ p7_a__8[31:23] ^ p7_a__8[8:0];
  assign p8_S0__92_comb = p7_a__8[11:2] ^ p7_a__8[22:13] ^ p7_a__8[31:22];
  assign p8_and_57219_comb = p7_a__8 & p7_a__7;
  assign p8_s_0__51_comb = p7_message[454:452] ^ p7_message[465:463];
  assign p8_s_0__50_comb = p7_message[451:448] ^ p7_message[462:459] ^ p7_message[479:476];
  assign p8_s_0__49_comb = p7_message[479:469] ^ p7_message[458:448] ^ p7_message[475:465];
  assign p8_s_0__48_comb = p7_message[468:455] ^ p7_message[479:466] ^ p7_message[464:451];
  assign p8_s_1__51_comb = p7_message[48:39] ^ p7_message[50:41];
  assign p8_s_1__50_comb = p7_message[38:32] ^ p7_message[40:34] ^ p7_message[63:57];
  assign p8_s_1__49_comb = p7_message[63:62] ^ p7_message[33:32] ^ p7_message[56:55];
  assign p8_s_1__48_comb = p7_message[61:49] ^ p7_message[63:51] ^ p7_message[54:42];
  assign p8_temp1__37_comb = p7_e__6 + p8_S1__9_comb;
  assign p8_ch__9_comb = p8_e__9_comb & p7_e__8 ^ ~(p8_e__9_comb | ~p7_e__7);
  assign p8_w_im15__8_comb = p7_message[223:192];
  assign p8_S0__8_comb = {p8_S0__95_comb, p8_S0__94_comb, p8_S0__93_comb, p8_S0__92_comb};
  assign p8_maj__8_comb = p8_and_57219_comb ^ p7_a__8 & p7_a__6 ^ p7_and_57141;
  assign p8_s_0__1_comb = {p8_s_0__51_comb, p8_s_0__50_comb, p8_s_0__49_comb, p8_s_0__48_comb};
  assign p8_s_1__1_comb = {p8_s_1__51_comb, p8_s_1__50_comb, p8_s_1__49_comb, p8_s_1__48_comb};
  assign p8_s_0__87_comb = p7_message[166:164] ^ p7_message[177:175];
  assign p8_s_0__86_comb = p7_message[163:160] ^ p7_message[174:171] ^ p7_message[191:188];
  assign p8_s_0__85_comb = p7_message[191:181] ^ p7_message[170:160] ^ p7_message[187:177];
  assign p8_s_0__84_comb = p7_message[180:167] ^ p7_message[191:178] ^ p7_message[176:163];
  assign p8_temp1__38_comb = p8_temp1__37_comb + p8_ch__9_comb;
  assign p8_temp1__267_comb = p8_w_im15__8_comb + 32'h1283_5b01;
  assign p8_temp2__8_comb = p8_S0__8_comb + p8_maj__8_comb;
  assign p8_value__1_comb = p7_message[511:480] + p8_s_0__1_comb;
  assign p8_value__2_comb = p8_w_im15__8_comb + p8_s_1__1_comb;
  assign p8_s_0__10_comb = {p8_s_0__87_comb, p8_s_0__86_comb, p8_s_0__85_comb, p8_s_0__84_comb};
  assign p8_temp1__40_comb = p8_temp1__38_comb + p8_temp1__267_comb;
  assign p8_a__9_comb = p7_temp1__436 + p8_temp2__8_comb;
  assign p8_value__3_comb = p8_value__1_comb + p8_value__2_comb;
  assign p8_value__28_comb = p8_w_im15__8_comb + p8_s_0__10_comb;

  // Registers for pipe stage 8:
  reg [511:0] p8_message;
  reg [31:0] p8_e__7;
  reg [31:0] p8_e__8;
  reg [31:0] p8_e__9;
  reg [31:0] p8_a__6;
  reg [31:0] p8_temp1__40;
  reg [31:0] p8_a__7;
  reg [31:0] p8_a__8;
  reg [31:0] p8_and_57219;
  reg [31:0] p8_a__9;
  reg [31:0] p8_value__3;
  reg [31:0] p8_value__7;
  reg [31:0] p8_value__13;
  reg [31:0] p8_value__16;
  reg [31:0] p8_value__22;
  reg [31:0] p8_value__28;
  always_ff @ (posedge clk) begin
    p8_message <= p7_message;
    p8_e__7 <= p7_e__7;
    p8_e__8 <= p7_e__8;
    p8_e__9 <= p8_e__9_comb;
    p8_a__6 <= p7_a__6;
    p8_temp1__40 <= p8_temp1__40_comb;
    p8_a__7 <= p7_a__7;
    p8_a__8 <= p7_a__8;
    p8_and_57219 <= p8_and_57219_comb;
    p8_a__9 <= p8_a__9_comb;
    p8_value__3 <= p8_value__3_comb;
    p8_value__7 <= p7_value__7;
    p8_value__13 <= p7_value__13;
    p8_value__16 <= p7_value__16;
    p8_value__22 <= p7_value__22;
    p8_value__28 <= p8_value__28_comb;
  end

  // ===== Pipe stage 9:
  wire [1:0] p9_S0__99_comb;
  wire [10:0] p9_S0__98_comb;
  wire [8:0] p9_S0__97_comb;
  wire [9:0] p9_S0__96_comb;
  wire [31:0] p9_and_57367_comb;
  wire [2:0] p9_s_0__55_comb;
  wire [3:0] p9_s_0__54_comb;
  wire [10:0] p9_s_0__53_comb;
  wire [13:0] p9_s_0__52_comb;
  wire [9:0] p9_s_1__55_comb;
  wire [6:0] p9_s_1__54_comb;
  wire [1:0] p9_s_1__53_comb;
  wire [12:0] p9_s_1__52_comb;
  wire [9:0] p9_s_1__59_comb;
  wire [6:0] p9_s_1__58_comb;
  wire [1:0] p9_s_1__57_comb;
  wire [12:0] p9_s_1__56_comb;
  wire [31:0] p9_S0__9_comb;
  wire [31:0] p9_maj__9_comb;
  wire [31:0] p9_w_init_im15_comb;
  wire [31:0] p9_s_0__2_comb;
  wire [31:0] p9_w_im15__9_comb;
  wire [31:0] p9_s_1__2_comb;
  wire [31:0] p9_w_im15__10_comb;
  wire [31:0] p9_s_1__3_comb;
  wire [31:0] p9_e__10_comb;
  wire [31:0] p9_temp2__9_comb;
  wire [31:0] p9_value__4_comb;
  wire [31:0] p9_value__5_comb;
  wire [31:0] p9_value__8_comb;
  wire [31:0] p9_a__10_comb;
  wire [31:0] p9_value__6_comb;
  wire [31:0] p9_value__9_comb;
  wire [5:0] p9_S1__103_comb;
  wire [4:0] p9_S1__102_comb;
  wire [13:0] p9_S1__101_comb;
  wire [6:0] p9_S1__100_comb;
  wire [30:0] p9_add_57332_comb;
  wire [31:0] p9_S1__10_comb;
  wire [31:0] p9_ch__10_comb;
  wire [31:0] p9_temp1__268_comb;
  wire [1:0] p9_S0__103_comb;
  wire [10:0] p9_S0__102_comb;
  wire [8:0] p9_S0__101_comb;
  wire [9:0] p9_S0__100_comb;
  wire [31:0] p9_and_57392_comb;
  wire [2:0] p9_s_0__63_comb;
  wire [3:0] p9_s_0__62_comb;
  wire [10:0] p9_s_0__61_comb;
  wire [13:0] p9_s_0__60_comb;
  wire [9:0] p9_s_1__63_comb;
  wire [6:0] p9_s_1__62_comb;
  wire [1:0] p9_s_1__61_comb;
  wire [12:0] p9_s_1__60_comb;
  wire [9:0] p9_s_1__67_comb;
  wire [6:0] p9_s_1__66_comb;
  wire [1:0] p9_s_1__65_comb;
  wire [12:0] p9_s_1__64_comb;
  wire [31:0] p9_temp1__431_comb;
  wire [31:0] p9_temp1__432_comb;
  wire [31:0] p9_S0__10_comb;
  wire [31:0] p9_maj__10_comb;
  wire [31:0] p9_w_im15__2_comb;
  wire [31:0] p9_s_0__4_comb;
  wire [31:0] p9_w_im15__11_comb;
  wire [31:0] p9_s_1__4_comb;
  wire [31:0] p9_w_im15__12_comb;
  wire [31:0] p9_s_1__5_comb;
  wire [2:0] p9_s_0__75_comb;
  wire [3:0] p9_s_0__74_comb;
  wire [10:0] p9_s_0__73_comb;
  wire [13:0] p9_s_0__72_comb;
  wire [2:0] p9_s_0__83_comb;
  wire [3:0] p9_s_0__82_comb;
  wire [10:0] p9_s_0__81_comb;
  wire [13:0] p9_s_0__80_comb;
  wire [2:0] p9_s_0__91_comb;
  wire [3:0] p9_s_0__90_comb;
  wire [10:0] p9_s_0__89_comb;
  wire [13:0] p9_s_0__88_comb;
  wire [2:0] p9_s_0__95_comb;
  wire [3:0] p9_s_0__94_comb;
  wire [10:0] p9_s_0__93_comb;
  wire [13:0] p9_s_0__92_comb;
  wire [2:0] p9_s_0__99_comb;
  wire [3:0] p9_s_0__98_comb;
  wire [10:0] p9_s_0__97_comb;
  wire [13:0] p9_s_0__96_comb;
  wire [2:0] p9_s_0__103_comb;
  wire [3:0] p9_s_0__102_comb;
  wire [10:0] p9_s_0__101_comb;
  wire [13:0] p9_s_0__100_comb;
  wire [2:0] p9_s_0__107_comb;
  wire [3:0] p9_s_0__106_comb;
  wire [10:0] p9_s_0__105_comb;
  wire [13:0] p9_s_0__104_comb;
  wire [31:0] p9_temp1__433_comb;
  wire [29:0] p9_add_57346_comb;
  wire [30:0] p9_add_57369_comb;
  wire [31:0] p9_temp2__10_comb;
  wire [29:0] p9_add_57401_comb;
  wire [31:0] p9_value__10_comb;
  wire [31:0] p9_value__11_comb;
  wire [31:0] p9_value__14_comb;
  wire [31:0] p9_w_im15__5_comb;
  wire [31:0] p9_s_0__7_comb;
  wire [31:0] p9_w_im15__7_comb;
  wire [31:0] p9_s_0__9_comb;
  wire [31:0] p9_s_0__11_comb;
  wire [31:0] p9_s_0__12_comb;
  wire [31:0] p9_s_0__13_comb;
  wire [31:0] p9_s_0__14_comb;
  wire [31:0] p9_w_init_im2_comb;
  wire [31:0] p9_s_0__15_comb;
  wire [31:0] p9_e__11_comb;
  wire [31:0] p9_temp1__269_comb;
  wire [31:0] p9_temp1__270_comb;
  wire [31:0] p9_temp1__271_comb;
  wire [31:0] p9_a__11_comb;
  wire [31:0] p9_temp1__273_comb;
  wire [31:0] p9_value__12_comb;
  wire [31:0] p9_value__15_comb;
  wire [31:0] p9_w_im2__1_comb;
  wire [31:0] p9_value__19_comb;
  wire [31:0] p9_value__25_comb;
  wire [31:0] p9_value__31_comb;
  wire [31:0] p9_value__34_comb;
  wire [31:0] p9_value__37_comb;
  wire [31:0] p9_value__40_comb;
  wire [31:0] p9_value__43_comb;
  assign p9_S0__99_comb = p8_a__9[1:0] ^ p8_a__9[12:11] ^ p8_a__9[21:20];
  assign p9_S0__98_comb = p8_a__9[31:21] ^ p8_a__9[10:0] ^ p8_a__9[19:9];
  assign p9_S0__97_comb = p8_a__9[20:12] ^ p8_a__9[31:23] ^ p8_a__9[8:0];
  assign p9_S0__96_comb = p8_a__9[11:2] ^ p8_a__9[22:13] ^ p8_a__9[31:22];
  assign p9_and_57367_comb = p8_a__9 & p8_a__8;
  assign p9_s_0__55_comb = p8_message[422:420] ^ p8_message[433:431];
  assign p9_s_0__54_comb = p8_message[419:416] ^ p8_message[430:427] ^ p8_message[447:444];
  assign p9_s_0__53_comb = p8_message[447:437] ^ p8_message[426:416] ^ p8_message[443:433];
  assign p9_s_0__52_comb = p8_message[436:423] ^ p8_message[447:434] ^ p8_message[432:419];
  assign p9_s_1__55_comb = p8_message[16:7] ^ p8_message[18:9];
  assign p9_s_1__54_comb = p8_message[6:0] ^ p8_message[8:2] ^ p8_message[31:25];
  assign p9_s_1__53_comb = p8_message[31:30] ^ p8_message[1:0] ^ p8_message[24:23];
  assign p9_s_1__52_comb = p8_message[29:17] ^ p8_message[31:19] ^ p8_message[22:10];
  assign p9_s_1__59_comb = p8_value__3[16:7] ^ p8_value__3[18:9];
  assign p9_s_1__58_comb = p8_value__3[6:0] ^ p8_value__3[8:2] ^ p8_value__3[31:25];
  assign p9_s_1__57_comb = p8_value__3[31:30] ^ p8_value__3[1:0] ^ p8_value__3[24:23];
  assign p9_s_1__56_comb = p8_value__3[29:17] ^ p8_value__3[31:19] ^ p8_value__3[22:10];
  assign p9_S0__9_comb = {p9_S0__99_comb, p9_S0__98_comb, p9_S0__97_comb, p9_S0__96_comb};
  assign p9_maj__9_comb = p9_and_57367_comb ^ p8_a__9 & p8_a__7 ^ p8_and_57219;
  assign p9_w_init_im15_comb = p8_message[479:448];
  assign p9_s_0__2_comb = {p9_s_0__55_comb, p9_s_0__54_comb, p9_s_0__53_comb, p9_s_0__52_comb};
  assign p9_w_im15__9_comb = p8_message[191:160];
  assign p9_s_1__2_comb = {p9_s_1__55_comb, p9_s_1__54_comb, p9_s_1__53_comb, p9_s_1__52_comb};
  assign p9_w_im15__10_comb = p8_message[159:128];
  assign p9_s_1__3_comb = {p9_s_1__59_comb, p9_s_1__58_comb, p9_s_1__57_comb, p9_s_1__56_comb};
  assign p9_e__10_comb = p8_a__6 + p8_temp1__40;
  assign p9_temp2__9_comb = p9_S0__9_comb + p9_maj__9_comb;
  assign p9_value__4_comb = p9_w_init_im15_comb + p9_s_0__2_comb;
  assign p9_value__5_comb = p9_w_im15__9_comb + p9_s_1__2_comb;
  assign p9_value__8_comb = p9_w_im15__10_comb + p9_s_1__3_comb;
  assign p9_a__10_comb = p8_temp1__40 + p9_temp2__9_comb;
  assign p9_value__6_comb = p9_value__4_comb + p9_value__5_comb;
  assign p9_value__9_comb = p8_value__7 + p9_value__8_comb;
  assign p9_S1__103_comb = p9_e__10_comb[5:0] ^ p9_e__10_comb[10:5] ^ p9_e__10_comb[24:19];
  assign p9_S1__102_comb = p9_e__10_comb[31:27] ^ p9_e__10_comb[4:0] ^ p9_e__10_comb[18:14];
  assign p9_S1__101_comb = p9_e__10_comb[26:13] ^ p9_e__10_comb[31:18] ^ p9_e__10_comb[13:0];
  assign p9_S1__100_comb = p9_e__10_comb[12:6] ^ p9_e__10_comb[17:11] ^ p9_e__10_comb[31:25];
  assign p9_add_57332_comb = p8_message[191:161] + 31'h1218_c2df;
  assign p9_S1__10_comb = {p9_S1__103_comb, p9_S1__102_comb, p9_S1__101_comb, p9_S1__100_comb};
  assign p9_ch__10_comb = p9_e__10_comb & p8_e__9 ^ ~(p9_e__10_comb | ~p8_e__8);
  assign p9_temp1__268_comb = {p9_add_57332_comb, p8_message[160]};
  assign p9_S0__103_comb = p9_a__10_comb[1:0] ^ p9_a__10_comb[12:11] ^ p9_a__10_comb[21:20];
  assign p9_S0__102_comb = p9_a__10_comb[31:21] ^ p9_a__10_comb[10:0] ^ p9_a__10_comb[19:9];
  assign p9_S0__101_comb = p9_a__10_comb[20:12] ^ p9_a__10_comb[31:23] ^ p9_a__10_comb[8:0];
  assign p9_S0__100_comb = p9_a__10_comb[11:2] ^ p9_a__10_comb[22:13] ^ p9_a__10_comb[31:22];
  assign p9_and_57392_comb = p9_a__10_comb & p8_a__9;
  assign p9_s_0__63_comb = p8_message[358:356] ^ p8_message[369:367];
  assign p9_s_0__62_comb = p8_message[355:352] ^ p8_message[366:363] ^ p8_message[383:380];
  assign p9_s_0__61_comb = p8_message[383:373] ^ p8_message[362:352] ^ p8_message[379:369];
  assign p9_s_0__60_comb = p8_message[372:359] ^ p8_message[383:370] ^ p8_message[368:355];
  assign p9_s_1__63_comb = p9_value__6_comb[16:7] ^ p9_value__6_comb[18:9];
  assign p9_s_1__62_comb = p9_value__6_comb[6:0] ^ p9_value__6_comb[8:2] ^ p9_value__6_comb[31:25];
  assign p9_s_1__61_comb = p9_value__6_comb[31:30] ^ p9_value__6_comb[1:0] ^ p9_value__6_comb[24:23];
  assign p9_s_1__60_comb = p9_value__6_comb[29:17] ^ p9_value__6_comb[31:19] ^ p9_value__6_comb[22:10];
  assign p9_s_1__67_comb = p9_value__9_comb[16:7] ^ p9_value__9_comb[18:9];
  assign p9_s_1__66_comb = p9_value__9_comb[6:0] ^ p9_value__9_comb[8:2] ^ p9_value__9_comb[31:25];
  assign p9_s_1__65_comb = p9_value__9_comb[31:30] ^ p9_value__9_comb[1:0] ^ p9_value__9_comb[24:23];
  assign p9_s_1__64_comb = p9_value__9_comb[29:17] ^ p9_value__9_comb[31:19] ^ p9_value__9_comb[22:10];
  assign p9_temp1__431_comb = p8_e__7 + p9_S1__10_comb;
  assign p9_temp1__432_comb = p9_ch__10_comb + p9_temp1__268_comb;
  assign p9_S0__10_comb = {p9_S0__103_comb, p9_S0__102_comb, p9_S0__101_comb, p9_S0__100_comb};
  assign p9_maj__10_comb = p9_and_57392_comb ^ p9_a__10_comb & p8_a__8 ^ p9_and_57367_comb;
  assign p9_w_im15__2_comb = p8_message[415:384];
  assign p9_s_0__4_comb = {p9_s_0__63_comb, p9_s_0__62_comb, p9_s_0__61_comb, p9_s_0__60_comb};
  assign p9_w_im15__11_comb = p8_message[127:96];
  assign p9_s_1__4_comb = {p9_s_1__63_comb, p9_s_1__62_comb, p9_s_1__61_comb, p9_s_1__60_comb};
  assign p9_w_im15__12_comb = p8_message[95:64];
  assign p9_s_1__5_comb = {p9_s_1__67_comb, p9_s_1__66_comb, p9_s_1__65_comb, p9_s_1__64_comb};
  assign p9_s_0__75_comb = p8_message[262:260] ^ p8_message[273:271];
  assign p9_s_0__74_comb = p8_message[259:256] ^ p8_message[270:267] ^ p8_message[287:284];
  assign p9_s_0__73_comb = p8_message[287:277] ^ p8_message[266:256] ^ p8_message[283:273];
  assign p9_s_0__72_comb = p8_message[276:263] ^ p8_message[287:274] ^ p8_message[272:259];
  assign p9_s_0__83_comb = p8_message[198:196] ^ p8_message[209:207];
  assign p9_s_0__82_comb = p8_message[195:192] ^ p8_message[206:203] ^ p8_message[223:220];
  assign p9_s_0__81_comb = p8_message[223:213] ^ p8_message[202:192] ^ p8_message[219:209];
  assign p9_s_0__80_comb = p8_message[212:199] ^ p8_message[223:210] ^ p8_message[208:195];
  assign p9_s_0__91_comb = p8_message[134:132] ^ p8_message[145:143];
  assign p9_s_0__90_comb = p8_message[131:128] ^ p8_message[142:139] ^ p8_message[159:156];
  assign p9_s_0__89_comb = p8_message[159:149] ^ p8_message[138:128] ^ p8_message[155:145];
  assign p9_s_0__88_comb = p8_message[148:135] ^ p8_message[159:146] ^ p8_message[144:131];
  assign p9_s_0__95_comb = p8_message[102:100] ^ p8_message[113:111];
  assign p9_s_0__94_comb = p8_message[99:96] ^ p8_message[110:107] ^ p8_message[127:124];
  assign p9_s_0__93_comb = p8_message[127:117] ^ p8_message[106:96] ^ p8_message[123:113];
  assign p9_s_0__92_comb = p8_message[116:103] ^ p8_message[127:114] ^ p8_message[112:99];
  assign p9_s_0__99_comb = p8_message[70:68] ^ p8_message[81:79];
  assign p9_s_0__98_comb = p8_message[67:64] ^ p8_message[78:75] ^ p8_message[95:92];
  assign p9_s_0__97_comb = p8_message[95:85] ^ p8_message[74:64] ^ p8_message[91:81];
  assign p9_s_0__96_comb = p8_message[84:71] ^ p8_message[95:82] ^ p8_message[80:67];
  assign p9_s_0__103_comb = p8_message[38:36] ^ p8_message[49:47];
  assign p9_s_0__102_comb = p8_message[35:32] ^ p8_message[46:43] ^ p8_message[63:60];
  assign p9_s_0__101_comb = p8_message[63:53] ^ p8_message[42:32] ^ p8_message[59:49];
  assign p9_s_0__100_comb = p8_message[52:39] ^ p8_message[63:50] ^ p8_message[48:35];
  assign p9_s_0__107_comb = p8_message[6:4] ^ p8_message[17:15];
  assign p9_s_0__106_comb = p8_message[3:0] ^ p8_message[14:11] ^ p8_message[31:28];
  assign p9_s_0__105_comb = p8_message[31:21] ^ p8_message[10:0] ^ p8_message[27:17];
  assign p9_s_0__104_comb = p8_message[20:7] ^ p8_message[31:18] ^ p8_message[16:3];
  assign p9_temp1__433_comb = p9_temp1__431_comb + p9_temp1__432_comb;
  assign p9_add_57346_comb = p8_message[127:98] + 30'h1caf_975d;
  assign p9_add_57369_comb = p8_message[95:65] + 31'h406f_58ff;
  assign p9_temp2__10_comb = p9_S0__10_comb + p9_maj__10_comb;
  assign p9_add_57401_comb = p8_message[31:2] + 30'h3066_fc5d;
  assign p9_value__10_comb = p9_w_im15__2_comb + p9_s_0__4_comb;
  assign p9_value__11_comb = p9_w_im15__11_comb + p9_s_1__4_comb;
  assign p9_value__14_comb = p9_w_im15__12_comb + p9_s_1__5_comb;
  assign p9_w_im15__5_comb = p8_message[319:288];
  assign p9_s_0__7_comb = {p9_s_0__75_comb, p9_s_0__74_comb, p9_s_0__73_comb, p9_s_0__72_comb};
  assign p9_w_im15__7_comb = p8_message[255:224];
  assign p9_s_0__9_comb = {p9_s_0__83_comb, p9_s_0__82_comb, p9_s_0__81_comb, p9_s_0__80_comb};
  assign p9_s_0__11_comb = {p9_s_0__91_comb, p9_s_0__90_comb, p9_s_0__89_comb, p9_s_0__88_comb};
  assign p9_s_0__12_comb = {p9_s_0__95_comb, p9_s_0__94_comb, p9_s_0__93_comb, p9_s_0__92_comb};
  assign p9_s_0__13_comb = {p9_s_0__99_comb, p9_s_0__98_comb, p9_s_0__97_comb, p9_s_0__96_comb};
  assign p9_s_0__14_comb = {p9_s_0__103_comb, p9_s_0__102_comb, p9_s_0__101_comb, p9_s_0__100_comb};
  assign p9_w_init_im2_comb = p8_message[63:32];
  assign p9_s_0__15_comb = {p9_s_0__107_comb, p9_s_0__106_comb, p9_s_0__105_comb, p9_s_0__104_comb};
  assign p9_e__11_comb = p8_a__7 + p9_temp1__433_comb;
  assign p9_temp1__269_comb = p9_w_im15__10_comb + 32'h550c_7dc3;
  assign p9_temp1__270_comb = {p9_add_57346_comb, p8_message[97:96]};
  assign p9_temp1__271_comb = {p9_add_57369_comb, p8_message[64]};
  assign p9_a__11_comb = p9_temp1__433_comb + p9_temp2__10_comb;
  assign p9_temp1__273_comb = {p9_add_57401_comb, p8_message[1:0]};
  assign p9_value__12_comb = p9_value__10_comb + p9_value__11_comb;
  assign p9_value__15_comb = p8_value__13 + p9_value__14_comb;
  assign p9_w_im2__1_comb = p8_message[31:0];
  assign p9_value__19_comb = p9_w_im15__5_comb + p9_s_0__7_comb;
  assign p9_value__25_comb = p9_w_im15__7_comb + p9_s_0__9_comb;
  assign p9_value__31_comb = p9_w_im15__9_comb + p9_s_0__11_comb;
  assign p9_value__34_comb = p9_w_im15__10_comb + p9_s_0__12_comb;
  assign p9_value__37_comb = p9_w_im15__11_comb + p9_s_0__13_comb;
  assign p9_value__40_comb = p9_w_im15__12_comb + p9_s_0__14_comb;
  assign p9_value__43_comb = p9_w_init_im2_comb + p9_s_0__15_comb;

  // Registers for pipe stage 9:
  reg [31:0] p9_e__8;
  reg [31:0] p9_e__9;
  reg [31:0] p9_e__10;
  reg [31:0] p9_e__11;
  reg [31:0] p9_temp1__269;
  reg [31:0] p9_a__8;
  reg [31:0] p9_temp1__270;
  reg [31:0] p9_a__9;
  reg [31:0] p9_temp1__271;
  reg [31:0] p9_a__10;
  reg [31:0] p9_and_57392;
  reg [31:0] p9_w_init_im2;
  reg [31:0] p9_a__11;
  reg [31:0] p9_temp1__273;
  reg [31:0] p9_value__3;
  reg [31:0] p9_value__6;
  reg [31:0] p9_value__9;
  reg [31:0] p9_value__12;
  reg [31:0] p9_value__15;
  reg [31:0] p9_value__16;
  reg [31:0] p9_w_im2__1;
  reg [31:0] p9_value__19;
  reg [31:0] p9_value__22;
  reg [31:0] p9_value__25;
  reg [31:0] p9_value__28;
  reg [31:0] p9_value__31;
  reg [31:0] p9_value__34;
  reg [31:0] p9_value__37;
  reg [31:0] p9_value__40;
  reg [31:0] p9_value__43;
  always_ff @ (posedge clk) begin
    p9_e__8 <= p8_e__8;
    p9_e__9 <= p8_e__9;
    p9_e__10 <= p9_e__10_comb;
    p9_e__11 <= p9_e__11_comb;
    p9_temp1__269 <= p9_temp1__269_comb;
    p9_a__8 <= p8_a__8;
    p9_temp1__270 <= p9_temp1__270_comb;
    p9_a__9 <= p8_a__9;
    p9_temp1__271 <= p9_temp1__271_comb;
    p9_a__10 <= p9_a__10_comb;
    p9_and_57392 <= p9_and_57392_comb;
    p9_w_init_im2 <= p9_w_init_im2_comb;
    p9_a__11 <= p9_a__11_comb;
    p9_temp1__273 <= p9_temp1__273_comb;
    p9_value__3 <= p8_value__3;
    p9_value__6 <= p9_value__6_comb;
    p9_value__9 <= p9_value__9_comb;
    p9_value__12 <= p9_value__12_comb;
    p9_value__15 <= p9_value__15_comb;
    p9_value__16 <= p8_value__16;
    p9_w_im2__1 <= p9_w_im2__1_comb;
    p9_value__19 <= p9_value__19_comb;
    p9_value__22 <= p8_value__22;
    p9_value__25 <= p9_value__25_comb;
    p9_value__28 <= p8_value__28;
    p9_value__31 <= p9_value__31_comb;
    p9_value__34 <= p9_value__34_comb;
    p9_value__37 <= p9_value__37_comb;
    p9_value__40 <= p9_value__40_comb;
    p9_value__43 <= p9_value__43_comb;
  end

  // ===== Pipe stage 10:
  wire [5:0] p10_S1__107_comb;
  wire [4:0] p10_S1__106_comb;
  wire [13:0] p10_S1__105_comb;
  wire [6:0] p10_S1__104_comb;
  wire [31:0] p10_S1__11_comb;
  wire [31:0] p10_temp1__45_comb;
  wire [31:0] p10_ch__11_comb;
  wire [1:0] p10_S0__107_comb;
  wire [10:0] p10_S0__106_comb;
  wire [8:0] p10_S0__105_comb;
  wire [9:0] p10_S0__104_comb;
  wire [31:0] p10_and_57737_comb;
  wire [9:0] p10_s_1__75_comb;
  wire [6:0] p10_s_1__74_comb;
  wire [1:0] p10_s_1__73_comb;
  wire [12:0] p10_s_1__72_comb;
  wire [31:0] p10_temp1__46_comb;
  wire [31:0] p10_S0__11_comb;
  wire [31:0] p10_maj__11_comb;
  wire [31:0] p10_s_1__7_comb;
  wire [2:0] p10_s_0__111_comb;
  wire [3:0] p10_s_0__110_comb;
  wire [10:0] p10_s_0__109_comb;
  wire [13:0] p10_s_0__108_comb;
  wire [31:0] p10_temp1__48_comb;
  wire [31:0] p10_temp2__11_comb;
  wire [31:0] p10_value__20_comb;
  wire [31:0] p10_s_0__16_comb;
  wire [31:0] p10_e__12_comb;
  wire [31:0] p10_a__12_comb;
  wire [31:0] p10_value__21_comb;
  wire [31:0] p10_value__46_comb;
  assign p10_S1__107_comb = p9_e__11[5:0] ^ p9_e__11[10:5] ^ p9_e__11[24:19];
  assign p10_S1__106_comb = p9_e__11[31:27] ^ p9_e__11[4:0] ^ p9_e__11[18:14];
  assign p10_S1__105_comb = p9_e__11[26:13] ^ p9_e__11[31:18] ^ p9_e__11[13:0];
  assign p10_S1__104_comb = p9_e__11[12:6] ^ p9_e__11[17:11] ^ p9_e__11[31:25];
  assign p10_S1__11_comb = {p10_S1__107_comb, p10_S1__106_comb, p10_S1__105_comb, p10_S1__104_comb};
  assign p10_temp1__45_comb = p9_e__8 + p10_S1__11_comb;
  assign p10_ch__11_comb = p9_e__11 & p9_e__10 ^ ~(p9_e__11 | ~p9_e__9);
  assign p10_S0__107_comb = p9_a__11[1:0] ^ p9_a__11[12:11] ^ p9_a__11[21:20];
  assign p10_S0__106_comb = p9_a__11[31:21] ^ p9_a__11[10:0] ^ p9_a__11[19:9];
  assign p10_S0__105_comb = p9_a__11[20:12] ^ p9_a__11[31:23] ^ p9_a__11[8:0];
  assign p10_S0__104_comb = p9_a__11[11:2] ^ p9_a__11[22:13] ^ p9_a__11[31:22];
  assign p10_and_57737_comb = p9_a__11 & p9_a__10;
  assign p10_s_1__75_comb = p9_value__15[16:7] ^ p9_value__15[18:9];
  assign p10_s_1__74_comb = p9_value__15[6:0] ^ p9_value__15[8:2] ^ p9_value__15[31:25];
  assign p10_s_1__73_comb = p9_value__15[31:30] ^ p9_value__15[1:0] ^ p9_value__15[24:23];
  assign p10_s_1__72_comb = p9_value__15[29:17] ^ p9_value__15[31:19] ^ p9_value__15[22:10];
  assign p10_temp1__46_comb = p10_temp1__45_comb + p10_ch__11_comb;
  assign p10_S0__11_comb = {p10_S0__107_comb, p10_S0__106_comb, p10_S0__105_comb, p10_S0__104_comb};
  assign p10_maj__11_comb = p10_and_57737_comb ^ p9_a__11 & p9_a__9 ^ p9_and_57392;
  assign p10_s_1__7_comb = {p10_s_1__75_comb, p10_s_1__74_comb, p10_s_1__73_comb, p10_s_1__72_comb};
  assign p10_s_0__111_comb = p9_value__3[6:4] ^ p9_value__3[17:15];
  assign p10_s_0__110_comb = p9_value__3[3:0] ^ p9_value__3[14:11] ^ p9_value__3[31:28];
  assign p10_s_0__109_comb = p9_value__3[31:21] ^ p9_value__3[10:0] ^ p9_value__3[27:17];
  assign p10_s_0__108_comb = p9_value__3[20:7] ^ p9_value__3[31:18] ^ p9_value__3[16:3];
  assign p10_temp1__48_comb = p10_temp1__46_comb + p9_temp1__269;
  assign p10_temp2__11_comb = p10_S0__11_comb + p10_maj__11_comb;
  assign p10_value__20_comb = p9_w_im2__1 + p10_s_1__7_comb;
  assign p10_s_0__16_comb = {p10_s_0__111_comb, p10_s_0__110_comb, p10_s_0__109_comb, p10_s_0__108_comb};
  assign p10_e__12_comb = p9_a__8 + p10_temp1__48_comb;
  assign p10_a__12_comb = p10_temp1__48_comb + p10_temp2__11_comb;
  assign p10_value__21_comb = p9_value__19 + p10_value__20_comb;
  assign p10_value__46_comb = p9_w_im2__1 + p10_s_0__16_comb;

  // Registers for pipe stage 10:
  reg [31:0] p10_e__9;
  reg [31:0] p10_e__10;
  reg [31:0] p10_e__11;
  reg [31:0] p10_e__12;
  reg [31:0] p10_temp1__270;
  reg [31:0] p10_a__9;
  reg [31:0] p10_temp1__271;
  reg [31:0] p10_a__10;
  reg [31:0] p10_w_init_im2;
  reg [31:0] p10_a__11;
  reg [31:0] p10_and_57737;
  reg [31:0] p10_temp1__273;
  reg [31:0] p10_a__12;
  reg [31:0] p10_value__3;
  reg [31:0] p10_value__6;
  reg [31:0] p10_value__9;
  reg [31:0] p10_value__12;
  reg [31:0] p10_value__15;
  reg [31:0] p10_value__16;
  reg [31:0] p10_value__21;
  reg [31:0] p10_value__22;
  reg [31:0] p10_value__25;
  reg [31:0] p10_value__28;
  reg [31:0] p10_value__31;
  reg [31:0] p10_value__34;
  reg [31:0] p10_value__37;
  reg [31:0] p10_value__40;
  reg [31:0] p10_value__43;
  reg [31:0] p10_value__46;
  always_ff @ (posedge clk) begin
    p10_e__9 <= p9_e__9;
    p10_e__10 <= p9_e__10;
    p10_e__11 <= p9_e__11;
    p10_e__12 <= p10_e__12_comb;
    p10_temp1__270 <= p9_temp1__270;
    p10_a__9 <= p9_a__9;
    p10_temp1__271 <= p9_temp1__271;
    p10_a__10 <= p9_a__10;
    p10_w_init_im2 <= p9_w_init_im2;
    p10_a__11 <= p9_a__11;
    p10_and_57737 <= p10_and_57737_comb;
    p10_temp1__273 <= p9_temp1__273;
    p10_a__12 <= p10_a__12_comb;
    p10_value__3 <= p9_value__3;
    p10_value__6 <= p9_value__6;
    p10_value__9 <= p9_value__9;
    p10_value__12 <= p9_value__12;
    p10_value__15 <= p9_value__15;
    p10_value__16 <= p9_value__16;
    p10_value__21 <= p10_value__21_comb;
    p10_value__22 <= p9_value__22;
    p10_value__25 <= p9_value__25;
    p10_value__28 <= p9_value__28;
    p10_value__31 <= p9_value__31;
    p10_value__34 <= p9_value__34;
    p10_value__37 <= p9_value__37;
    p10_value__40 <= p9_value__40;
    p10_value__43 <= p9_value__43;
    p10_value__46 <= p10_value__46_comb;
  end

  // ===== Pipe stage 11:
  wire [5:0] p11_S1__111_comb;
  wire [4:0] p11_S1__110_comb;
  wire [13:0] p11_S1__109_comb;
  wire [6:0] p11_S1__108_comb;
  wire [31:0] p11_S1__12_comb;
  wire [31:0] p11_ch__12_comb;
  wire [31:0] p11_temp1__428_comb;
  wire [31:0] p11_temp1__429_comb;
  wire [31:0] p11_temp1__430_comb;
  wire [31:0] p11_e__13_comb;
  wire [1:0] p11_S0__111_comb;
  wire [10:0] p11_S0__110_comb;
  wire [8:0] p11_S0__109_comb;
  wire [9:0] p11_S0__108_comb;
  wire [31:0] p11_and_57900_comb;
  wire [5:0] p11_S1__115_comb;
  wire [4:0] p11_S1__114_comb;
  wire [13:0] p11_S1__113_comb;
  wire [6:0] p11_S1__112_comb;
  wire [31:0] p11_S0__12_comb;
  wire [31:0] p11_maj__12_comb;
  wire [31:0] p11_S1__13_comb;
  wire [31:0] p11_ch__13_comb;
  wire [31:0] p11_temp2__12_comb;
  wire [31:0] p11_temp1__425_comb;
  wire [31:0] p11_temp1__426_comb;
  wire [31:0] p11_a__13_comb;
  assign p11_S1__111_comb = p10_e__12[5:0] ^ p10_e__12[10:5] ^ p10_e__12[24:19];
  assign p11_S1__110_comb = p10_e__12[31:27] ^ p10_e__12[4:0] ^ p10_e__12[18:14];
  assign p11_S1__109_comb = p10_e__12[26:13] ^ p10_e__12[31:18] ^ p10_e__12[13:0];
  assign p11_S1__108_comb = p10_e__12[12:6] ^ p10_e__12[17:11] ^ p10_e__12[31:25];
  assign p11_S1__12_comb = {p11_S1__111_comb, p11_S1__110_comb, p11_S1__109_comb, p11_S1__108_comb};
  assign p11_ch__12_comb = p10_e__12 & p10_e__11 ^ ~(p10_e__12 | ~p10_e__10);
  assign p11_temp1__428_comb = p10_e__9 + p11_S1__12_comb;
  assign p11_temp1__429_comb = p11_ch__12_comb + p10_temp1__270;
  assign p11_temp1__430_comb = p11_temp1__428_comb + p11_temp1__429_comb;
  assign p11_e__13_comb = p10_a__9 + p11_temp1__430_comb;
  assign p11_S0__111_comb = p10_a__12[1:0] ^ p10_a__12[12:11] ^ p10_a__12[21:20];
  assign p11_S0__110_comb = p10_a__12[31:21] ^ p10_a__12[10:0] ^ p10_a__12[19:9];
  assign p11_S0__109_comb = p10_a__12[20:12] ^ p10_a__12[31:23] ^ p10_a__12[8:0];
  assign p11_S0__108_comb = p10_a__12[11:2] ^ p10_a__12[22:13] ^ p10_a__12[31:22];
  assign p11_and_57900_comb = p10_a__12 & p10_a__11;
  assign p11_S1__115_comb = p11_e__13_comb[5:0] ^ p11_e__13_comb[10:5] ^ p11_e__13_comb[24:19];
  assign p11_S1__114_comb = p11_e__13_comb[31:27] ^ p11_e__13_comb[4:0] ^ p11_e__13_comb[18:14];
  assign p11_S1__113_comb = p11_e__13_comb[26:13] ^ p11_e__13_comb[31:18] ^ p11_e__13_comb[13:0];
  assign p11_S1__112_comb = p11_e__13_comb[12:6] ^ p11_e__13_comb[17:11] ^ p11_e__13_comb[31:25];
  assign p11_S0__12_comb = {p11_S0__111_comb, p11_S0__110_comb, p11_S0__109_comb, p11_S0__108_comb};
  assign p11_maj__12_comb = p11_and_57900_comb ^ p10_a__12 & p10_a__10 ^ p10_and_57737;
  assign p11_S1__13_comb = {p11_S1__115_comb, p11_S1__114_comb, p11_S1__113_comb, p11_S1__112_comb};
  assign p11_ch__13_comb = p11_e__13_comb & p10_e__12 ^ ~(p11_e__13_comb | ~p10_e__11);
  assign p11_temp2__12_comb = p11_S0__12_comb + p11_maj__12_comb;
  assign p11_temp1__425_comb = p10_e__10 + p11_S1__13_comb;
  assign p11_temp1__426_comb = p11_ch__13_comb + p10_temp1__271;
  assign p11_a__13_comb = p11_temp1__430_comb + p11_temp2__12_comb;

  // Registers for pipe stage 11:
  reg [31:0] p11_e__11;
  reg [31:0] p11_e__12;
  reg [31:0] p11_e__13;
  reg [31:0] p11_temp1__425;
  reg [31:0] p11_temp1__426;
  reg [31:0] p11_a__10;
  reg [31:0] p11_w_init_im2;
  reg [31:0] p11_a__11;
  reg [31:0] p11_temp1__273;
  reg [31:0] p11_a__12;
  reg [31:0] p11_and_57900;
  reg [31:0] p11_value__3;
  reg [31:0] p11_a__13;
  reg [31:0] p11_value__6;
  reg [31:0] p11_value__9;
  reg [31:0] p11_value__12;
  reg [31:0] p11_value__15;
  reg [31:0] p11_value__16;
  reg [31:0] p11_value__21;
  reg [31:0] p11_value__22;
  reg [31:0] p11_value__25;
  reg [31:0] p11_value__28;
  reg [31:0] p11_value__31;
  reg [31:0] p11_value__34;
  reg [31:0] p11_value__37;
  reg [31:0] p11_value__40;
  reg [31:0] p11_value__43;
  reg [31:0] p11_value__46;
  always_ff @ (posedge clk) begin
    p11_e__11 <= p10_e__11;
    p11_e__12 <= p10_e__12;
    p11_e__13 <= p11_e__13_comb;
    p11_temp1__425 <= p11_temp1__425_comb;
    p11_temp1__426 <= p11_temp1__426_comb;
    p11_a__10 <= p10_a__10;
    p11_w_init_im2 <= p10_w_init_im2;
    p11_a__11 <= p10_a__11;
    p11_temp1__273 <= p10_temp1__273;
    p11_a__12 <= p10_a__12;
    p11_and_57900 <= p11_and_57900_comb;
    p11_value__3 <= p10_value__3;
    p11_a__13 <= p11_a__13_comb;
    p11_value__6 <= p10_value__6;
    p11_value__9 <= p10_value__9;
    p11_value__12 <= p10_value__12;
    p11_value__15 <= p10_value__15;
    p11_value__16 <= p10_value__16;
    p11_value__21 <= p10_value__21;
    p11_value__22 <= p10_value__22;
    p11_value__25 <= p10_value__25;
    p11_value__28 <= p10_value__28;
    p11_value__31 <= p10_value__31;
    p11_value__34 <= p10_value__34;
    p11_value__37 <= p10_value__37;
    p11_value__40 <= p10_value__40;
    p11_value__43 <= p10_value__43;
    p11_value__46 <= p10_value__46;
  end

  // ===== Pipe stage 12:
  wire [1:0] p12_bit_slice_58011_comb;
  wire [9:0] p12_s_1__71_comb;
  wire [6:0] p12_s_1__70_comb;
  wire [1:0] p12_s_1__69_comb;
  wire [12:0] p12_s_1__68_comb;
  wire [31:0] p12_s_1__6_comb;
  wire [31:0] p12_temp1__427_comb;
  wire [31:0] p12_value__17_comb;
  wire [31:0] p12_e__14_comb;
  wire [31:0] p12_value__18_comb;
  wire [5:0] p12_S1__119_comb;
  wire [4:0] p12_S1__118_comb;
  wire [13:0] p12_S1__117_comb;
  wire [6:0] p12_S1__116_comb;
  wire [1:0] p12_S0__115_comb;
  wire [10:0] p12_S0__114_comb;
  wire [8:0] p12_S0__113_comb;
  wire [9:0] p12_S0__112_comb;
  wire [31:0] p12_and_58005_comb;
  wire [9:0] p12_s_1__79_comb;
  wire [6:0] p12_s_1__78_comb;
  wire [1:0] p12_s_1__77_comb;
  wire [12:0] p12_s_1__76_comb;
  wire [31:0] p12_S1__14_comb;
  wire [31:0] p12_S0__13_comb;
  wire [31:0] p12_maj__13_comb;
  wire [31:0] p12_s_1__8_comb;
  wire [31:0] p12_temp1__57_comb;
  wire [31:0] p12_ch__14_comb;
  wire [31:0] p12_temp2__13_comb;
  wire [31:0] p12_value__23_comb;
  wire [31:0] p12_temp1__58_comb;
  wire [31:0] p12_temp1__272_comb;
  wire [31:0] p12_a__14_comb;
  wire [31:0] p12_value__24_comb;
  assign p12_bit_slice_58011_comb = p11_value__12[1:0];
  assign p12_s_1__71_comb = p11_value__12[16:7] ^ p11_value__12[18:9];
  assign p12_s_1__70_comb = p11_value__12[6:0] ^ p11_value__12[8:2] ^ p11_value__12[31:25];
  assign p12_s_1__69_comb = p11_value__12[31:30] ^ p12_bit_slice_58011_comb ^ p11_value__12[24:23];
  assign p12_s_1__68_comb = p11_value__12[29:17] ^ p11_value__12[31:19] ^ p11_value__12[22:10];
  assign p12_s_1__6_comb = {p12_s_1__71_comb, p12_s_1__70_comb, p12_s_1__69_comb, p12_s_1__68_comb};
  assign p12_temp1__427_comb = p11_temp1__425 + p11_temp1__426;
  assign p12_value__17_comb = p11_w_init_im2 + p12_s_1__6_comb;
  assign p12_e__14_comb = p11_a__10 + p12_temp1__427_comb;
  assign p12_value__18_comb = p11_value__16 + p12_value__17_comb;
  assign p12_S1__119_comb = p12_e__14_comb[5:0] ^ p12_e__14_comb[10:5] ^ p12_e__14_comb[24:19];
  assign p12_S1__118_comb = p12_e__14_comb[31:27] ^ p12_e__14_comb[4:0] ^ p12_e__14_comb[18:14];
  assign p12_S1__117_comb = p12_e__14_comb[26:13] ^ p12_e__14_comb[31:18] ^ p12_e__14_comb[13:0];
  assign p12_S1__116_comb = p12_e__14_comb[12:6] ^ p12_e__14_comb[17:11] ^ p12_e__14_comb[31:25];
  assign p12_S0__115_comb = p11_a__13[1:0] ^ p11_a__13[12:11] ^ p11_a__13[21:20];
  assign p12_S0__114_comb = p11_a__13[31:21] ^ p11_a__13[10:0] ^ p11_a__13[19:9];
  assign p12_S0__113_comb = p11_a__13[20:12] ^ p11_a__13[31:23] ^ p11_a__13[8:0];
  assign p12_S0__112_comb = p11_a__13[11:2] ^ p11_a__13[22:13] ^ p11_a__13[31:22];
  assign p12_and_58005_comb = p11_a__13 & p11_a__12;
  assign p12_s_1__79_comb = p12_value__18_comb[16:7] ^ p12_value__18_comb[18:9];
  assign p12_s_1__78_comb = p12_value__18_comb[6:0] ^ p12_value__18_comb[8:2] ^ p12_value__18_comb[31:25];
  assign p12_s_1__77_comb = p12_value__18_comb[31:30] ^ p12_value__18_comb[1:0] ^ p12_value__18_comb[24:23];
  assign p12_s_1__76_comb = p12_value__18_comb[29:17] ^ p12_value__18_comb[31:19] ^ p12_value__18_comb[22:10];
  assign p12_S1__14_comb = {p12_S1__119_comb, p12_S1__118_comb, p12_S1__117_comb, p12_S1__116_comb};
  assign p12_S0__13_comb = {p12_S0__115_comb, p12_S0__114_comb, p12_S0__113_comb, p12_S0__112_comb};
  assign p12_maj__13_comb = p12_and_58005_comb ^ p11_a__13 & p11_a__11 ^ p11_and_57900;
  assign p12_s_1__8_comb = {p12_s_1__79_comb, p12_s_1__78_comb, p12_s_1__77_comb, p12_s_1__76_comb};
  assign p12_temp1__57_comb = p11_e__11 + p12_S1__14_comb;
  assign p12_ch__14_comb = p12_e__14_comb & p11_e__13 ^ ~(p12_e__14_comb | ~p11_e__12);
  assign p12_temp2__13_comb = p12_S0__13_comb + p12_maj__13_comb;
  assign p12_value__23_comb = p11_value__3 + p12_s_1__8_comb;
  assign p12_temp1__58_comb = p12_temp1__57_comb + p12_ch__14_comb;
  assign p12_temp1__272_comb = p11_w_init_im2 + 32'h9bdc_06a7;
  assign p12_a__14_comb = p12_temp1__427_comb + p12_temp2__13_comb;
  assign p12_value__24_comb = p11_value__22 + p12_value__23_comb;

  // Registers for pipe stage 12:
  reg [31:0] p12_e__12;
  reg [31:0] p12_e__13;
  reg [31:0] p12_e__14;
  reg [31:0] p12_temp1__58;
  reg [31:0] p12_temp1__272;
  reg [31:0] p12_a__11;
  reg [31:0] p12_temp1__273;
  reg [31:0] p12_a__12;
  reg [31:0] p12_value__3;
  reg [31:0] p12_a__13;
  reg [31:0] p12_value__6;
  reg [31:0] p12_and_58005;
  reg [31:0] p12_a__14;
  reg [31:0] p12_value__9;
  reg [31:0] p12_value__12;
  reg [1:0] p12_bit_slice_58011;
  reg [31:0] p12_value__15;
  reg [31:0] p12_value__18;
  reg [31:0] p12_value__21;
  reg [31:0] p12_value__24;
  reg [31:0] p12_value__25;
  reg [31:0] p12_value__28;
  reg [31:0] p12_value__31;
  reg [31:0] p12_value__34;
  reg [31:0] p12_value__37;
  reg [31:0] p12_value__40;
  reg [31:0] p12_value__43;
  reg [31:0] p12_value__46;
  always_ff @ (posedge clk) begin
    p12_e__12 <= p11_e__12;
    p12_e__13 <= p11_e__13;
    p12_e__14 <= p12_e__14_comb;
    p12_temp1__58 <= p12_temp1__58_comb;
    p12_temp1__272 <= p12_temp1__272_comb;
    p12_a__11 <= p11_a__11;
    p12_temp1__273 <= p11_temp1__273;
    p12_a__12 <= p11_a__12;
    p12_value__3 <= p11_value__3;
    p12_a__13 <= p11_a__13;
    p12_value__6 <= p11_value__6;
    p12_and_58005 <= p12_and_58005_comb;
    p12_a__14 <= p12_a__14_comb;
    p12_value__9 <= p11_value__9;
    p12_value__12 <= p11_value__12;
    p12_bit_slice_58011 <= p12_bit_slice_58011_comb;
    p12_value__15 <= p11_value__15;
    p12_value__18 <= p12_value__18_comb;
    p12_value__21 <= p11_value__21;
    p12_value__24 <= p12_value__24_comb;
    p12_value__25 <= p11_value__25;
    p12_value__28 <= p11_value__28;
    p12_value__31 <= p11_value__31;
    p12_value__34 <= p11_value__34;
    p12_value__37 <= p11_value__37;
    p12_value__40 <= p11_value__40;
    p12_value__43 <= p11_value__43;
    p12_value__46 <= p11_value__46;
  end

  // ===== Pipe stage 13:
  wire [9:0] p13_s_1__87_comb;
  wire [6:0] p13_s_1__86_comb;
  wire [1:0] p13_s_1__85_comb;
  wire [12:0] p13_s_1__84_comb;
  wire [31:0] p13_s_1__10_comb;
  wire [31:0] p13_temp1__60_comb;
  wire [31:0] p13_value__29_comb;
  wire [31:0] p13_e__15_comb;
  wire [31:0] p13_value__30_comb;
  wire [5:0] p13_S1__123_comb;
  wire [4:0] p13_S1__122_comb;
  wire [13:0] p13_S1__121_comb;
  wire [6:0] p13_S1__120_comb;
  wire [1:0] p13_S0__119_comb;
  wire [10:0] p13_S0__118_comb;
  wire [8:0] p13_S0__117_comb;
  wire [9:0] p13_S0__116_comb;
  wire [31:0] p13_and_58145_comb;
  wire [9:0] p13_s_1__95_comb;
  wire [6:0] p13_s_1__94_comb;
  wire [1:0] p13_s_1__93_comb;
  wire [12:0] p13_s_1__92_comb;
  wire [31:0] p13_S1__15_comb;
  wire [31:0] p13_ch__15_comb;
  wire [31:0] p13_S0__14_comb;
  wire [31:0] p13_maj__14_comb;
  wire [31:0] p13_s_1__12_comb;
  wire [31:0] p13_temp1__422_comb;
  wire [31:0] p13_temp1__423_comb;
  wire [31:0] p13_temp2__14_comb;
  wire [31:0] p13_value__35_comb;
  wire [31:0] p13_temp1__424_comb;
  wire [31:0] p13_a__15_comb;
  wire [31:0] p13_value__36_comb;
  assign p13_s_1__87_comb = p12_value__24[16:7] ^ p12_value__24[18:9];
  assign p13_s_1__86_comb = p12_value__24[6:0] ^ p12_value__24[8:2] ^ p12_value__24[31:25];
  assign p13_s_1__85_comb = p12_value__24[31:30] ^ p12_value__24[1:0] ^ p12_value__24[24:23];
  assign p13_s_1__84_comb = p12_value__24[29:17] ^ p12_value__24[31:19] ^ p12_value__24[22:10];
  assign p13_s_1__10_comb = {p13_s_1__87_comb, p13_s_1__86_comb, p13_s_1__85_comb, p13_s_1__84_comb};
  assign p13_temp1__60_comb = p12_temp1__58 + p12_temp1__272;
  assign p13_value__29_comb = p12_value__9 + p13_s_1__10_comb;
  assign p13_e__15_comb = p12_a__11 + p13_temp1__60_comb;
  assign p13_value__30_comb = p12_value__28 + p13_value__29_comb;
  assign p13_S1__123_comb = p13_e__15_comb[5:0] ^ p13_e__15_comb[10:5] ^ p13_e__15_comb[24:19];
  assign p13_S1__122_comb = p13_e__15_comb[31:27] ^ p13_e__15_comb[4:0] ^ p13_e__15_comb[18:14];
  assign p13_S1__121_comb = p13_e__15_comb[26:13] ^ p13_e__15_comb[31:18] ^ p13_e__15_comb[13:0];
  assign p13_S1__120_comb = p13_e__15_comb[12:6] ^ p13_e__15_comb[17:11] ^ p13_e__15_comb[31:25];
  assign p13_S0__119_comb = p12_a__14[1:0] ^ p12_a__14[12:11] ^ p12_a__14[21:20];
  assign p13_S0__118_comb = p12_a__14[31:21] ^ p12_a__14[10:0] ^ p12_a__14[19:9];
  assign p13_S0__117_comb = p12_a__14[20:12] ^ p12_a__14[31:23] ^ p12_a__14[8:0];
  assign p13_S0__116_comb = p12_a__14[11:2] ^ p12_a__14[22:13] ^ p12_a__14[31:22];
  assign p13_and_58145_comb = p12_a__14 & p12_a__13;
  assign p13_s_1__95_comb = p13_value__30_comb[16:7] ^ p13_value__30_comb[18:9];
  assign p13_s_1__94_comb = p13_value__30_comb[6:0] ^ p13_value__30_comb[8:2] ^ p13_value__30_comb[31:25];
  assign p13_s_1__93_comb = p13_value__30_comb[31:30] ^ p13_value__30_comb[1:0] ^ p13_value__30_comb[24:23];
  assign p13_s_1__92_comb = p13_value__30_comb[29:17] ^ p13_value__30_comb[31:19] ^ p13_value__30_comb[22:10];
  assign p13_S1__15_comb = {p13_S1__123_comb, p13_S1__122_comb, p13_S1__121_comb, p13_S1__120_comb};
  assign p13_ch__15_comb = p13_e__15_comb & p12_e__14 ^ ~(p13_e__15_comb | ~p12_e__13);
  assign p13_S0__14_comb = {p13_S0__119_comb, p13_S0__118_comb, p13_S0__117_comb, p13_S0__116_comb};
  assign p13_maj__14_comb = p13_and_58145_comb ^ p12_a__14 & p12_a__12 ^ p12_and_58005;
  assign p13_s_1__12_comb = {p13_s_1__95_comb, p13_s_1__94_comb, p13_s_1__93_comb, p13_s_1__92_comb};
  assign p13_temp1__422_comb = p12_e__12 + p13_S1__15_comb;
  assign p13_temp1__423_comb = p13_ch__15_comb + p12_temp1__273;
  assign p13_temp2__14_comb = p13_S0__14_comb + p13_maj__14_comb;
  assign p13_value__35_comb = p12_value__15 + p13_s_1__12_comb;
  assign p13_temp1__424_comb = p13_temp1__422_comb + p13_temp1__423_comb;
  assign p13_a__15_comb = p13_temp1__60_comb + p13_temp2__14_comb;
  assign p13_value__36_comb = p12_value__34 + p13_value__35_comb;

  // Registers for pipe stage 13:
  reg [31:0] p13_e__13;
  reg [31:0] p13_e__14;
  reg [31:0] p13_e__15;
  reg [31:0] p13_a__12;
  reg [31:0] p13_temp1__424;
  reg [31:0] p13_value__3;
  reg [31:0] p13_a__13;
  reg [31:0] p13_value__6;
  reg [31:0] p13_a__14;
  reg [31:0] p13_value__9;
  reg [31:0] p13_and_58145;
  reg [31:0] p13_a__15;
  reg [31:0] p13_value__12;
  reg [1:0] p13_bit_slice_58011;
  reg [31:0] p13_value__15;
  reg [31:0] p13_value__18;
  reg [31:0] p13_value__21;
  reg [31:0] p13_value__24;
  reg [31:0] p13_value__25;
  reg [31:0] p13_value__30;
  reg [31:0] p13_value__31;
  reg [31:0] p13_value__36;
  reg [31:0] p13_value__37;
  reg [31:0] p13_value__40;
  reg [31:0] p13_value__43;
  reg [31:0] p13_value__46;
  always_ff @ (posedge clk) begin
    p13_e__13 <= p12_e__13;
    p13_e__14 <= p12_e__14;
    p13_e__15 <= p13_e__15_comb;
    p13_a__12 <= p12_a__12;
    p13_temp1__424 <= p13_temp1__424_comb;
    p13_value__3 <= p12_value__3;
    p13_a__13 <= p12_a__13;
    p13_value__6 <= p12_value__6;
    p13_a__14 <= p12_a__14;
    p13_value__9 <= p12_value__9;
    p13_and_58145 <= p13_and_58145_comb;
    p13_a__15 <= p13_a__15_comb;
    p13_value__12 <= p12_value__12;
    p13_bit_slice_58011 <= p12_bit_slice_58011;
    p13_value__15 <= p12_value__15;
    p13_value__18 <= p12_value__18;
    p13_value__21 <= p12_value__21;
    p13_value__24 <= p12_value__24;
    p13_value__25 <= p12_value__25;
    p13_value__30 <= p13_value__30_comb;
    p13_value__31 <= p12_value__31;
    p13_value__36 <= p13_value__36_comb;
    p13_value__37 <= p12_value__37;
    p13_value__40 <= p12_value__40;
    p13_value__43 <= p12_value__43;
    p13_value__46 <= p12_value__46;
  end

  // ===== Pipe stage 14:
  wire [31:0] p14_e__16_comb;
  wire [5:0] p14_S1__127_comb;
  wire [4:0] p14_S1__126_comb;
  wire [13:0] p14_S1__125_comb;
  wire [6:0] p14_S1__124_comb;
  wire [31:0] p14_S1__16_comb;
  wire [1:0] p14_S0__123_comb;
  wire [10:0] p14_S0__122_comb;
  wire [8:0] p14_S0__121_comb;
  wire [9:0] p14_S0__120_comb;
  wire [31:0] p14_and_58282_comb;
  wire [9:0] p14_s_1__103_comb;
  wire [6:0] p14_s_1__102_comb;
  wire [1:0] p14_s_1__101_comb;
  wire [12:0] p14_s_1__100_comb;
  wire [31:0] p14_temp1__65_comb;
  wire [31:0] p14_ch__16_comb;
  wire [31:0] p14_S0__15_comb;
  wire [31:0] p14_maj__15_comb;
  wire [31:0] p14_s_1__14_comb;
  wire [2:0] p14_s_0__115_comb;
  wire [3:0] p14_s_0__114_comb;
  wire [10:0] p14_s_0__113_comb;
  wire [13:0] p14_s_0__112_comb;
  wire [31:0] p14_temp1__66_comb;
  wire [31:0] p14_temp1__274_comb;
  wire [31:0] p14_temp2__15_comb;
  wire [31:0] p14_value__41_comb;
  wire [31:0] p14_s_0__17_comb;
  wire [31:0] p14_temp1__68_comb;
  wire [31:0] p14_a__16_comb;
  wire [31:0] p14_value__42_comb;
  wire [31:0] p14_value__49_comb;
  assign p14_e__16_comb = p13_a__12 + p13_temp1__424;
  assign p14_S1__127_comb = p14_e__16_comb[5:0] ^ p14_e__16_comb[10:5] ^ p14_e__16_comb[24:19];
  assign p14_S1__126_comb = p14_e__16_comb[31:27] ^ p14_e__16_comb[4:0] ^ p14_e__16_comb[18:14];
  assign p14_S1__125_comb = p14_e__16_comb[26:13] ^ p14_e__16_comb[31:18] ^ p14_e__16_comb[13:0];
  assign p14_S1__124_comb = p14_e__16_comb[12:6] ^ p14_e__16_comb[17:11] ^ p14_e__16_comb[31:25];
  assign p14_S1__16_comb = {p14_S1__127_comb, p14_S1__126_comb, p14_S1__125_comb, p14_S1__124_comb};
  assign p14_S0__123_comb = p13_a__15[1:0] ^ p13_a__15[12:11] ^ p13_a__15[21:20];
  assign p14_S0__122_comb = p13_a__15[31:21] ^ p13_a__15[10:0] ^ p13_a__15[19:9];
  assign p14_S0__121_comb = p13_a__15[20:12] ^ p13_a__15[31:23] ^ p13_a__15[8:0];
  assign p14_S0__120_comb = p13_a__15[11:2] ^ p13_a__15[22:13] ^ p13_a__15[31:22];
  assign p14_and_58282_comb = p13_a__15 & p13_a__14;
  assign p14_s_1__103_comb = p13_value__36[16:7] ^ p13_value__36[18:9];
  assign p14_s_1__102_comb = p13_value__36[6:0] ^ p13_value__36[8:2] ^ p13_value__36[31:25];
  assign p14_s_1__101_comb = p13_value__36[31:30] ^ p13_value__36[1:0] ^ p13_value__36[24:23];
  assign p14_s_1__100_comb = p13_value__36[29:17] ^ p13_value__36[31:19] ^ p13_value__36[22:10];
  assign p14_temp1__65_comb = p13_e__13 + p14_S1__16_comb;
  assign p14_ch__16_comb = p14_e__16_comb & p13_e__15 ^ ~(p14_e__16_comb | ~p13_e__14);
  assign p14_S0__15_comb = {p14_S0__123_comb, p14_S0__122_comb, p14_S0__121_comb, p14_S0__120_comb};
  assign p14_maj__15_comb = p14_and_58282_comb ^ p13_a__15 & p13_a__13 ^ p13_and_58145;
  assign p14_s_1__14_comb = {p14_s_1__103_comb, p14_s_1__102_comb, p14_s_1__101_comb, p14_s_1__100_comb};
  assign p14_s_0__115_comb = p13_value__6[6:4] ^ p13_value__6[17:15];
  assign p14_s_0__114_comb = p13_value__6[3:0] ^ p13_value__6[14:11] ^ p13_value__6[31:28];
  assign p14_s_0__113_comb = p13_value__6[31:21] ^ p13_value__6[10:0] ^ p13_value__6[27:17];
  assign p14_s_0__112_comb = p13_value__6[20:7] ^ p13_value__6[31:18] ^ p13_value__6[16:3];
  assign p14_temp1__66_comb = p14_temp1__65_comb + p14_ch__16_comb;
  assign p14_temp1__274_comb = p13_value__3 + 32'he49b_69c1;
  assign p14_temp2__15_comb = p14_S0__15_comb + p14_maj__15_comb;
  assign p14_value__41_comb = p13_value__21 + p14_s_1__14_comb;
  assign p14_s_0__17_comb = {p14_s_0__115_comb, p14_s_0__114_comb, p14_s_0__113_comb, p14_s_0__112_comb};
  assign p14_temp1__68_comb = p14_temp1__66_comb + p14_temp1__274_comb;
  assign p14_a__16_comb = p13_temp1__424 + p14_temp2__15_comb;
  assign p14_value__42_comb = p13_value__40 + p14_value__41_comb;
  assign p14_value__49_comb = p13_value__3 + p14_s_0__17_comb;

  // Registers for pipe stage 14:
  reg [31:0] p14_e__14;
  reg [31:0] p14_e__15;
  reg [31:0] p14_e__16;
  reg [31:0] p14_a__13;
  reg [31:0] p14_temp1__68;
  reg [31:0] p14_value__6;
  reg [31:0] p14_a__14;
  reg [31:0] p14_value__9;
  reg [31:0] p14_a__15;
  reg [31:0] p14_value__12;
  reg [31:0] p14_and_58282;
  reg [1:0] p14_bit_slice_58011;
  reg [31:0] p14_a__16;
  reg [31:0] p14_value__15;
  reg [31:0] p14_value__18;
  reg [31:0] p14_value__21;
  reg [31:0] p14_value__24;
  reg [31:0] p14_value__25;
  reg [31:0] p14_value__30;
  reg [31:0] p14_value__31;
  reg [31:0] p14_value__36;
  reg [31:0] p14_value__37;
  reg [31:0] p14_value__42;
  reg [31:0] p14_value__43;
  reg [31:0] p14_value__46;
  reg [31:0] p14_value__49;
  always_ff @ (posedge clk) begin
    p14_e__14 <= p13_e__14;
    p14_e__15 <= p13_e__15;
    p14_e__16 <= p14_e__16_comb;
    p14_a__13 <= p13_a__13;
    p14_temp1__68 <= p14_temp1__68_comb;
    p14_value__6 <= p13_value__6;
    p14_a__14 <= p13_a__14;
    p14_value__9 <= p13_value__9;
    p14_a__15 <= p13_a__15;
    p14_value__12 <= p13_value__12;
    p14_and_58282 <= p14_and_58282_comb;
    p14_bit_slice_58011 <= p13_bit_slice_58011;
    p14_a__16 <= p14_a__16_comb;
    p14_value__15 <= p13_value__15;
    p14_value__18 <= p13_value__18;
    p14_value__21 <= p13_value__21;
    p14_value__24 <= p13_value__24;
    p14_value__25 <= p13_value__25;
    p14_value__30 <= p13_value__30;
    p14_value__31 <= p13_value__31;
    p14_value__36 <= p13_value__36;
    p14_value__37 <= p13_value__37;
    p14_value__42 <= p14_value__42_comb;
    p14_value__43 <= p13_value__43;
    p14_value__46 <= p13_value__46;
    p14_value__49 <= p14_value__49_comb;
  end

  // ===== Pipe stage 15:
  wire [1:0] p15_S0__127_comb;
  wire [10:0] p15_S0__126_comb;
  wire [8:0] p15_S0__125_comb;
  wire [9:0] p15_S0__124_comb;
  wire [31:0] p15_and_58425_comb;
  wire [31:0] p15_S0__16_comb;
  wire [31:0] p15_maj__16_comb;
  wire [31:0] p15_e__17_comb;
  wire [31:0] p15_temp2__16_comb;
  wire [31:0] p15_a__17_comb;
  wire [5:0] p15_S1__131_comb;
  wire [4:0] p15_S1__130_comb;
  wire [13:0] p15_S1__129_comb;
  wire [6:0] p15_S1__128_comb;
  wire [30:0] p15_add_58397_comb;
  wire [31:0] p15_S1__17_comb;
  wire [31:0] p15_ch__17_comb;
  wire [31:0] p15_temp1__275_comb;
  wire [1:0] p15_S0__131_comb;
  wire [10:0] p15_S0__130_comb;
  wire [8:0] p15_S0__129_comb;
  wire [9:0] p15_S0__128_comb;
  wire [31:0] p15_and_58447_comb;
  wire [31:0] p15_temp1__419_comb;
  wire [31:0] p15_temp1__420_comb;
  wire [31:0] p15_S0__17_comb;
  wire [31:0] p15_maj__17_comb;
  wire [31:0] p15_temp1__421_comb;
  wire [31:0] p15_temp2__17_comb;
  wire [31:0] p15_e__18_comb;
  wire [30:0] p15_add_58408_comb;
  wire [31:0] p15_a__18_comb;
  assign p15_S0__127_comb = p14_a__16[1:0] ^ p14_a__16[12:11] ^ p14_a__16[21:20];
  assign p15_S0__126_comb = p14_a__16[31:21] ^ p14_a__16[10:0] ^ p14_a__16[19:9];
  assign p15_S0__125_comb = p14_a__16[20:12] ^ p14_a__16[31:23] ^ p14_a__16[8:0];
  assign p15_S0__124_comb = p14_a__16[11:2] ^ p14_a__16[22:13] ^ p14_a__16[31:22];
  assign p15_and_58425_comb = p14_a__16 & p14_a__15;
  assign p15_S0__16_comb = {p15_S0__127_comb, p15_S0__126_comb, p15_S0__125_comb, p15_S0__124_comb};
  assign p15_maj__16_comb = p15_and_58425_comb ^ p14_a__16 & p14_a__14 ^ p14_and_58282;
  assign p15_e__17_comb = p14_a__13 + p14_temp1__68;
  assign p15_temp2__16_comb = p15_S0__16_comb + p15_maj__16_comb;
  assign p15_a__17_comb = p14_temp1__68 + p15_temp2__16_comb;
  assign p15_S1__131_comb = p15_e__17_comb[5:0] ^ p15_e__17_comb[10:5] ^ p15_e__17_comb[24:19];
  assign p15_S1__130_comb = p15_e__17_comb[31:27] ^ p15_e__17_comb[4:0] ^ p15_e__17_comb[18:14];
  assign p15_S1__129_comb = p15_e__17_comb[26:13] ^ p15_e__17_comb[31:18] ^ p15_e__17_comb[13:0];
  assign p15_S1__128_comb = p15_e__17_comb[12:6] ^ p15_e__17_comb[17:11] ^ p15_e__17_comb[31:25];
  assign p15_add_58397_comb = p14_value__6[31:1] + 31'h77df_23c3;
  assign p15_S1__17_comb = {p15_S1__131_comb, p15_S1__130_comb, p15_S1__129_comb, p15_S1__128_comb};
  assign p15_ch__17_comb = p15_e__17_comb & p14_e__16 ^ ~(p15_e__17_comb | ~p14_e__15);
  assign p15_temp1__275_comb = {p15_add_58397_comb, p14_value__6[0]};
  assign p15_S0__131_comb = p15_a__17_comb[1:0] ^ p15_a__17_comb[12:11] ^ p15_a__17_comb[21:20];
  assign p15_S0__130_comb = p15_a__17_comb[31:21] ^ p15_a__17_comb[10:0] ^ p15_a__17_comb[19:9];
  assign p15_S0__129_comb = p15_a__17_comb[20:12] ^ p15_a__17_comb[31:23] ^ p15_a__17_comb[8:0];
  assign p15_S0__128_comb = p15_a__17_comb[11:2] ^ p15_a__17_comb[22:13] ^ p15_a__17_comb[31:22];
  assign p15_and_58447_comb = p15_a__17_comb & p14_a__16;
  assign p15_temp1__419_comb = p14_e__14 + p15_S1__17_comb;
  assign p15_temp1__420_comb = p15_ch__17_comb + p15_temp1__275_comb;
  assign p15_S0__17_comb = {p15_S0__131_comb, p15_S0__130_comb, p15_S0__129_comb, p15_S0__128_comb};
  assign p15_maj__17_comb = p15_and_58447_comb ^ p15_a__17_comb & p14_a__15 ^ p15_and_58425_comb;
  assign p15_temp1__421_comb = p15_temp1__419_comb + p15_temp1__420_comb;
  assign p15_temp2__17_comb = p15_S0__17_comb + p15_maj__17_comb;
  assign p15_e__18_comb = p14_a__14 + p15_temp1__421_comb;
  assign p15_add_58408_comb = p14_value__9[31:1] + 31'h07e0_cee3;
  assign p15_a__18_comb = p15_temp1__421_comb + p15_temp2__17_comb;

  // Registers for pipe stage 15:
  reg [31:0] p15_e__15;
  reg [31:0] p15_e__16;
  reg [31:0] p15_e__17;
  reg [31:0] p15_value__6;
  reg [31:0] p15_e__18;
  reg [31:0] p15_value__9;
  reg [30:0] p15_add_58408;
  reg [31:0] p15_a__15;
  reg [31:0] p15_value__12;
  reg [1:0] p15_bit_slice_58011;
  reg [31:0] p15_a__16;
  reg [31:0] p15_value__15;
  reg [31:0] p15_a__17;
  reg [31:0] p15_value__18;
  reg [31:0] p15_and_58447;
  reg [31:0] p15_a__18;
  reg [31:0] p15_value__21;
  reg [31:0] p15_value__24;
  reg [31:0] p15_value__25;
  reg [31:0] p15_value__30;
  reg [31:0] p15_value__31;
  reg [31:0] p15_value__36;
  reg [31:0] p15_value__37;
  reg [31:0] p15_value__42;
  reg [31:0] p15_value__43;
  reg [31:0] p15_value__46;
  reg [31:0] p15_value__49;
  always_ff @ (posedge clk) begin
    p15_e__15 <= p14_e__15;
    p15_e__16 <= p14_e__16;
    p15_e__17 <= p15_e__17_comb;
    p15_value__6 <= p14_value__6;
    p15_e__18 <= p15_e__18_comb;
    p15_value__9 <= p14_value__9;
    p15_add_58408 <= p15_add_58408_comb;
    p15_a__15 <= p14_a__15;
    p15_value__12 <= p14_value__12;
    p15_bit_slice_58011 <= p14_bit_slice_58011;
    p15_a__16 <= p14_a__16;
    p15_value__15 <= p14_value__15;
    p15_a__17 <= p15_a__17_comb;
    p15_value__18 <= p14_value__18;
    p15_and_58447 <= p15_and_58447_comb;
    p15_a__18 <= p15_a__18_comb;
    p15_value__21 <= p14_value__21;
    p15_value__24 <= p14_value__24;
    p15_value__25 <= p14_value__25;
    p15_value__30 <= p14_value__30;
    p15_value__31 <= p14_value__31;
    p15_value__36 <= p14_value__36;
    p15_value__37 <= p14_value__37;
    p15_value__42 <= p14_value__42;
    p15_value__43 <= p14_value__43;
    p15_value__46 <= p14_value__46;
    p15_value__49 <= p14_value__49;
  end

  // ===== Pipe stage 16:
  wire [5:0] p16_S1__135_comb;
  wire [4:0] p16_S1__134_comb;
  wire [13:0] p16_S1__133_comb;
  wire [6:0] p16_S1__132_comb;
  wire [31:0] p16_S1__18_comb;
  wire [31:0] p16_ch__18_comb;
  wire [31:0] p16_temp1__276_comb;
  wire [31:0] p16_temp1__416_comb;
  wire [31:0] p16_temp1__417_comb;
  wire [31:0] p16_temp1__418_comb;
  wire [31:0] p16_e__19_comb;
  wire [1:0] p16_S0__135_comb;
  wire [10:0] p16_S0__134_comb;
  wire [8:0] p16_S0__133_comb;
  wire [9:0] p16_S0__132_comb;
  wire [31:0] p16_and_58577_comb;
  wire [5:0] p16_S1__139_comb;
  wire [4:0] p16_S1__138_comb;
  wire [13:0] p16_S1__137_comb;
  wire [6:0] p16_S1__136_comb;
  wire [29:0] p16_add_58555_comb;
  wire [31:0] p16_S0__18_comb;
  wire [31:0] p16_maj__18_comb;
  wire [31:0] p16_S1__19_comb;
  wire [31:0] p16_ch__19_comb;
  wire [31:0] p16_temp1__277_comb;
  wire [31:0] p16_temp2__18_comb;
  wire [31:0] p16_temp1__413_comb;
  wire [31:0] p16_temp1__414_comb;
  wire [31:0] p16_a__19_comb;
  assign p16_S1__135_comb = p15_e__18[5:0] ^ p15_e__18[10:5] ^ p15_e__18[24:19];
  assign p16_S1__134_comb = p15_e__18[31:27] ^ p15_e__18[4:0] ^ p15_e__18[18:14];
  assign p16_S1__133_comb = p15_e__18[26:13] ^ p15_e__18[31:18] ^ p15_e__18[13:0];
  assign p16_S1__132_comb = p15_e__18[12:6] ^ p15_e__18[17:11] ^ p15_e__18[31:25];
  assign p16_S1__18_comb = {p16_S1__135_comb, p16_S1__134_comb, p16_S1__133_comb, p16_S1__132_comb};
  assign p16_ch__18_comb = p15_e__18 & p15_e__17 ^ ~(p15_e__18 | ~p15_e__16);
  assign p16_temp1__276_comb = {p15_add_58408, p15_value__9[0]};
  assign p16_temp1__416_comb = p15_e__15 + p16_S1__18_comb;
  assign p16_temp1__417_comb = p16_ch__18_comb + p16_temp1__276_comb;
  assign p16_temp1__418_comb = p16_temp1__416_comb + p16_temp1__417_comb;
  assign p16_e__19_comb = p15_a__15 + p16_temp1__418_comb;
  assign p16_S0__135_comb = p15_a__18[1:0] ^ p15_a__18[12:11] ^ p15_a__18[21:20];
  assign p16_S0__134_comb = p15_a__18[31:21] ^ p15_a__18[10:0] ^ p15_a__18[19:9];
  assign p16_S0__133_comb = p15_a__18[20:12] ^ p15_a__18[31:23] ^ p15_a__18[8:0];
  assign p16_S0__132_comb = p15_a__18[11:2] ^ p15_a__18[22:13] ^ p15_a__18[31:22];
  assign p16_and_58577_comb = p15_a__18 & p15_a__17;
  assign p16_S1__139_comb = p16_e__19_comb[5:0] ^ p16_e__19_comb[10:5] ^ p16_e__19_comb[24:19];
  assign p16_S1__138_comb = p16_e__19_comb[31:27] ^ p16_e__19_comb[4:0] ^ p16_e__19_comb[18:14];
  assign p16_S1__137_comb = p16_e__19_comb[26:13] ^ p16_e__19_comb[31:18] ^ p16_e__19_comb[13:0];
  assign p16_S1__136_comb = p16_e__19_comb[12:6] ^ p16_e__19_comb[17:11] ^ p16_e__19_comb[31:25];
  assign p16_add_58555_comb = p15_value__12[31:2] + 30'h0903_2873;
  assign p16_S0__18_comb = {p16_S0__135_comb, p16_S0__134_comb, p16_S0__133_comb, p16_S0__132_comb};
  assign p16_maj__18_comb = p16_and_58577_comb ^ p15_a__18 & p15_a__16 ^ p15_and_58447;
  assign p16_S1__19_comb = {p16_S1__139_comb, p16_S1__138_comb, p16_S1__137_comb, p16_S1__136_comb};
  assign p16_ch__19_comb = p16_e__19_comb & p15_e__18 ^ ~(p16_e__19_comb | ~p15_e__17);
  assign p16_temp1__277_comb = {p16_add_58555_comb, p15_bit_slice_58011};
  assign p16_temp2__18_comb = p16_S0__18_comb + p16_maj__18_comb;
  assign p16_temp1__413_comb = p15_e__16 + p16_S1__19_comb;
  assign p16_temp1__414_comb = p16_ch__19_comb + p16_temp1__277_comb;
  assign p16_a__19_comb = p16_temp1__418_comb + p16_temp2__18_comb;

  // Registers for pipe stage 16:
  reg [31:0] p16_e__17;
  reg [31:0] p16_value__6;
  reg [31:0] p16_e__18;
  reg [31:0] p16_value__9;
  reg [31:0] p16_e__19;
  reg [31:0] p16_value__12;
  reg [31:0] p16_temp1__413;
  reg [31:0] p16_temp1__414;
  reg [31:0] p16_a__16;
  reg [31:0] p16_value__15;
  reg [31:0] p16_a__17;
  reg [31:0] p16_value__18;
  reg [31:0] p16_a__18;
  reg [31:0] p16_value__21;
  reg [31:0] p16_and_58577;
  reg [31:0] p16_a__19;
  reg [31:0] p16_value__24;
  reg [31:0] p16_value__25;
  reg [31:0] p16_value__30;
  reg [31:0] p16_value__31;
  reg [31:0] p16_value__36;
  reg [31:0] p16_value__37;
  reg [31:0] p16_value__42;
  reg [31:0] p16_value__43;
  reg [31:0] p16_value__46;
  reg [31:0] p16_value__49;
  always_ff @ (posedge clk) begin
    p16_e__17 <= p15_e__17;
    p16_value__6 <= p15_value__6;
    p16_e__18 <= p15_e__18;
    p16_value__9 <= p15_value__9;
    p16_e__19 <= p16_e__19_comb;
    p16_value__12 <= p15_value__12;
    p16_temp1__413 <= p16_temp1__413_comb;
    p16_temp1__414 <= p16_temp1__414_comb;
    p16_a__16 <= p15_a__16;
    p16_value__15 <= p15_value__15;
    p16_a__17 <= p15_a__17;
    p16_value__18 <= p15_value__18;
    p16_a__18 <= p15_a__18;
    p16_value__21 <= p15_value__21;
    p16_and_58577 <= p16_and_58577_comb;
    p16_a__19 <= p16_a__19_comb;
    p16_value__24 <= p15_value__24;
    p16_value__25 <= p15_value__25;
    p16_value__30 <= p15_value__30;
    p16_value__31 <= p15_value__31;
    p16_value__36 <= p15_value__36;
    p16_value__37 <= p15_value__37;
    p16_value__42 <= p15_value__42;
    p16_value__43 <= p15_value__43;
    p16_value__46 <= p15_value__46;
    p16_value__49 <= p15_value__49;
  end

  // ===== Pipe stage 17:
  wire [31:0] p17_temp1__415_comb;
  wire [31:0] p17_e__20_comb;
  wire [5:0] p17_S1__143_comb;
  wire [4:0] p17_S1__142_comb;
  wire [13:0] p17_S1__141_comb;
  wire [6:0] p17_S1__140_comb;
  wire [1:0] p17_S0__139_comb;
  wire [10:0] p17_S0__138_comb;
  wire [8:0] p17_S0__137_comb;
  wire [9:0] p17_S0__136_comb;
  wire [31:0] p17_and_58678_comb;
  wire [31:0] p17_S1__20_comb;
  wire [31:0] p17_S0__19_comb;
  wire [31:0] p17_maj__19_comb;
  wire [31:0] p17_temp1__81_comb;
  wire [31:0] p17_ch__20_comb;
  wire [31:0] p17_temp2__19_comb;
  wire [31:0] p17_temp1__82_comb;
  wire [31:0] p17_temp1__278_comb;
  wire [31:0] p17_a__20_comb;
  assign p17_temp1__415_comb = p16_temp1__413 + p16_temp1__414;
  assign p17_e__20_comb = p16_a__16 + p17_temp1__415_comb;
  assign p17_S1__143_comb = p17_e__20_comb[5:0] ^ p17_e__20_comb[10:5] ^ p17_e__20_comb[24:19];
  assign p17_S1__142_comb = p17_e__20_comb[31:27] ^ p17_e__20_comb[4:0] ^ p17_e__20_comb[18:14];
  assign p17_S1__141_comb = p17_e__20_comb[26:13] ^ p17_e__20_comb[31:18] ^ p17_e__20_comb[13:0];
  assign p17_S1__140_comb = p17_e__20_comb[12:6] ^ p17_e__20_comb[17:11] ^ p17_e__20_comb[31:25];
  assign p17_S0__139_comb = p16_a__19[1:0] ^ p16_a__19[12:11] ^ p16_a__19[21:20];
  assign p17_S0__138_comb = p16_a__19[31:21] ^ p16_a__19[10:0] ^ p16_a__19[19:9];
  assign p17_S0__137_comb = p16_a__19[20:12] ^ p16_a__19[31:23] ^ p16_a__19[8:0];
  assign p17_S0__136_comb = p16_a__19[11:2] ^ p16_a__19[22:13] ^ p16_a__19[31:22];
  assign p17_and_58678_comb = p16_a__19 & p16_a__18;
  assign p17_S1__20_comb = {p17_S1__143_comb, p17_S1__142_comb, p17_S1__141_comb, p17_S1__140_comb};
  assign p17_S0__19_comb = {p17_S0__139_comb, p17_S0__138_comb, p17_S0__137_comb, p17_S0__136_comb};
  assign p17_maj__19_comb = p17_and_58678_comb ^ p16_a__19 & p16_a__17 ^ p16_and_58577;
  assign p17_temp1__81_comb = p16_e__17 + p17_S1__20_comb;
  assign p17_ch__20_comb = p17_e__20_comb & p16_e__19 ^ ~(p17_e__20_comb | ~p16_e__18);
  assign p17_temp2__19_comb = p17_S0__19_comb + p17_maj__19_comb;
  assign p17_temp1__82_comb = p17_temp1__81_comb + p17_ch__20_comb;
  assign p17_temp1__278_comb = p16_value__15 + 32'h2de9_2c6f;
  assign p17_a__20_comb = p17_temp1__415_comb + p17_temp2__19_comb;

  // Registers for pipe stage 17:
  reg [31:0] p17_value__6;
  reg [31:0] p17_e__18;
  reg [31:0] p17_value__9;
  reg [31:0] p17_e__19;
  reg [31:0] p17_value__12;
  reg [31:0] p17_e__20;
  reg [31:0] p17_value__15;
  reg [31:0] p17_temp1__82;
  reg [31:0] p17_temp1__278;
  reg [31:0] p17_a__17;
  reg [31:0] p17_value__18;
  reg [31:0] p17_a__18;
  reg [31:0] p17_value__21;
  reg [31:0] p17_a__19;
  reg [31:0] p17_value__24;
  reg [31:0] p17_and_58678;
  reg [31:0] p17_a__20;
  reg [31:0] p17_value__25;
  reg [31:0] p17_value__30;
  reg [31:0] p17_value__31;
  reg [31:0] p17_value__36;
  reg [31:0] p17_value__37;
  reg [31:0] p17_value__42;
  reg [31:0] p17_value__43;
  reg [31:0] p17_value__46;
  reg [31:0] p17_value__49;
  always_ff @ (posedge clk) begin
    p17_value__6 <= p16_value__6;
    p17_e__18 <= p16_e__18;
    p17_value__9 <= p16_value__9;
    p17_e__19 <= p16_e__19;
    p17_value__12 <= p16_value__12;
    p17_e__20 <= p17_e__20_comb;
    p17_value__15 <= p16_value__15;
    p17_temp1__82 <= p17_temp1__82_comb;
    p17_temp1__278 <= p17_temp1__278_comb;
    p17_a__17 <= p16_a__17;
    p17_value__18 <= p16_value__18;
    p17_a__18 <= p16_a__18;
    p17_value__21 <= p16_value__21;
    p17_a__19 <= p16_a__19;
    p17_value__24 <= p16_value__24;
    p17_and_58678 <= p17_and_58678_comb;
    p17_a__20 <= p17_a__20_comb;
    p17_value__25 <= p16_value__25;
    p17_value__30 <= p16_value__30;
    p17_value__31 <= p16_value__31;
    p17_value__36 <= p16_value__36;
    p17_value__37 <= p16_value__37;
    p17_value__42 <= p16_value__42;
    p17_value__43 <= p16_value__43;
    p17_value__46 <= p16_value__46;
    p17_value__49 <= p16_value__49;
  end

  // ===== Pipe stage 18:
  wire [31:0] p18_temp1__84_comb;
  wire [31:0] p18_e__21_comb;
  wire [5:0] p18_S1__147_comb;
  wire [4:0] p18_S1__146_comb;
  wire [13:0] p18_S1__145_comb;
  wire [6:0] p18_S1__144_comb;
  wire [30:0] p18_add_58759_comb;
  wire [1:0] p18_S0__143_comb;
  wire [10:0] p18_S0__142_comb;
  wire [8:0] p18_S0__141_comb;
  wire [9:0] p18_S0__140_comb;
  wire [31:0] p18_and_58783_comb;
  wire [31:0] p18_S1__21_comb;
  wire [31:0] p18_ch__21_comb;
  wire [31:0] p18_temp1__279_comb;
  wire [31:0] p18_S0__20_comb;
  wire [31:0] p18_maj__20_comb;
  wire [31:0] p18_temp1__410_comb;
  wire [31:0] p18_temp1__411_comb;
  wire [31:0] p18_temp2__20_comb;
  wire [31:0] p18_temp1__412_comb;
  wire [31:0] p18_a__21_comb;
  assign p18_temp1__84_comb = p17_temp1__82 + p17_temp1__278;
  assign p18_e__21_comb = p17_a__17 + p18_temp1__84_comb;
  assign p18_S1__147_comb = p18_e__21_comb[5:0] ^ p18_e__21_comb[10:5] ^ p18_e__21_comb[24:19];
  assign p18_S1__146_comb = p18_e__21_comb[31:27] ^ p18_e__21_comb[4:0] ^ p18_e__21_comb[18:14];
  assign p18_S1__145_comb = p18_e__21_comb[26:13] ^ p18_e__21_comb[31:18] ^ p18_e__21_comb[13:0];
  assign p18_S1__144_comb = p18_e__21_comb[12:6] ^ p18_e__21_comb[17:11] ^ p18_e__21_comb[31:25];
  assign p18_add_58759_comb = p17_value__18[31:1] + 31'h253a_4255;
  assign p18_S0__143_comb = p17_a__20[1:0] ^ p17_a__20[12:11] ^ p17_a__20[21:20];
  assign p18_S0__142_comb = p17_a__20[31:21] ^ p17_a__20[10:0] ^ p17_a__20[19:9];
  assign p18_S0__141_comb = p17_a__20[20:12] ^ p17_a__20[31:23] ^ p17_a__20[8:0];
  assign p18_S0__140_comb = p17_a__20[11:2] ^ p17_a__20[22:13] ^ p17_a__20[31:22];
  assign p18_and_58783_comb = p17_a__20 & p17_a__19;
  assign p18_S1__21_comb = {p18_S1__147_comb, p18_S1__146_comb, p18_S1__145_comb, p18_S1__144_comb};
  assign p18_ch__21_comb = p18_e__21_comb & p17_e__20 ^ ~(p18_e__21_comb | ~p17_e__19);
  assign p18_temp1__279_comb = {p18_add_58759_comb, p17_value__18[0]};
  assign p18_S0__20_comb = {p18_S0__143_comb, p18_S0__142_comb, p18_S0__141_comb, p18_S0__140_comb};
  assign p18_maj__20_comb = p18_and_58783_comb ^ p17_a__20 & p17_a__18 ^ p17_and_58678;
  assign p18_temp1__410_comb = p17_e__18 + p18_S1__21_comb;
  assign p18_temp1__411_comb = p18_ch__21_comb + p18_temp1__279_comb;
  assign p18_temp2__20_comb = p18_S0__20_comb + p18_maj__20_comb;
  assign p18_temp1__412_comb = p18_temp1__410_comb + p18_temp1__411_comb;
  assign p18_a__21_comb = p18_temp1__84_comb + p18_temp2__20_comb;

  // Registers for pipe stage 18:
  reg [31:0] p18_value__6;
  reg [31:0] p18_value__9;
  reg [31:0] p18_e__19;
  reg [31:0] p18_value__12;
  reg [31:0] p18_e__20;
  reg [31:0] p18_value__15;
  reg [31:0] p18_e__21;
  reg [31:0] p18_value__18;
  reg [31:0] p18_a__18;
  reg [31:0] p18_temp1__412;
  reg [31:0] p18_value__21;
  reg [31:0] p18_a__19;
  reg [31:0] p18_value__24;
  reg [31:0] p18_a__20;
  reg [31:0] p18_value__25;
  reg [31:0] p18_and_58783;
  reg [31:0] p18_a__21;
  reg [31:0] p18_value__30;
  reg [31:0] p18_value__31;
  reg [31:0] p18_value__36;
  reg [31:0] p18_value__37;
  reg [31:0] p18_value__42;
  reg [31:0] p18_value__43;
  reg [31:0] p18_value__46;
  reg [31:0] p18_value__49;
  always_ff @ (posedge clk) begin
    p18_value__6 <= p17_value__6;
    p18_value__9 <= p17_value__9;
    p18_e__19 <= p17_e__19;
    p18_value__12 <= p17_value__12;
    p18_e__20 <= p17_e__20;
    p18_value__15 <= p17_value__15;
    p18_e__21 <= p18_e__21_comb;
    p18_value__18 <= p17_value__18;
    p18_a__18 <= p17_a__18;
    p18_temp1__412 <= p18_temp1__412_comb;
    p18_value__21 <= p17_value__21;
    p18_a__19 <= p17_a__19;
    p18_value__24 <= p17_value__24;
    p18_a__20 <= p17_a__20;
    p18_value__25 <= p17_value__25;
    p18_and_58783 <= p18_and_58783_comb;
    p18_a__21 <= p18_a__21_comb;
    p18_value__30 <= p17_value__30;
    p18_value__31 <= p17_value__31;
    p18_value__36 <= p17_value__36;
    p18_value__37 <= p17_value__37;
    p18_value__42 <= p17_value__42;
    p18_value__43 <= p17_value__43;
    p18_value__46 <= p17_value__46;
    p18_value__49 <= p17_value__49;
  end

  // ===== Pipe stage 19:
  wire [9:0] p19_s_1__83_comb;
  wire [6:0] p19_s_1__82_comb;
  wire [1:0] p19_s_1__81_comb;
  wire [12:0] p19_s_1__80_comb;
  wire [1:0] p19_S0__147_comb;
  wire [10:0] p19_S0__146_comb;
  wire [8:0] p19_S0__145_comb;
  wire [9:0] p19_S0__144_comb;
  wire [31:0] p19_and_58906_comb;
  wire [31:0] p19_s_1__9_comb;
  wire [31:0] p19_S0__21_comb;
  wire [31:0] p19_maj__21_comb;
  wire [31:0] p19_e__22_comb;
  wire [31:0] p19_value__26_comb;
  wire [31:0] p19_temp2__21_comb;
  wire [31:0] p19_value__27_comb;
  wire [31:0] p19_a__22_comb;
  wire [5:0] p19_S1__151_comb;
  wire [4:0] p19_S1__150_comb;
  wire [13:0] p19_S1__149_comb;
  wire [6:0] p19_S1__148_comb;
  wire [29:0] p19_add_58861_comb;
  wire [31:0] p19_S1__22_comb;
  wire [31:0] p19_ch__22_comb;
  wire [31:0] p19_temp1__280_comb;
  wire [9:0] p19_s_1__91_comb;
  wire [6:0] p19_s_1__90_comb;
  wire [1:0] p19_s_1__89_comb;
  wire [12:0] p19_s_1__88_comb;
  wire [1:0] p19_S0__151_comb;
  wire [10:0] p19_S0__150_comb;
  wire [8:0] p19_S0__149_comb;
  wire [9:0] p19_S0__148_comb;
  wire [31:0] p19_and_58946_comb;
  wire [9:0] p19_s_1__111_comb;
  wire [6:0] p19_s_1__110_comb;
  wire [1:0] p19_s_1__109_comb;
  wire [12:0] p19_s_1__108_comb;
  wire [31:0] p19_temp1__407_comb;
  wire [31:0] p19_temp1__408_comb;
  wire [31:0] p19_s_1__11_comb;
  wire [31:0] p19_S0__22_comb;
  wire [31:0] p19_maj__22_comb;
  wire [31:0] p19_s_1__16_comb;
  wire [2:0] p19_s_0__119_comb;
  wire [3:0] p19_s_0__118_comb;
  wire [10:0] p19_s_0__117_comb;
  wire [13:0] p19_s_0__116_comb;
  wire [2:0] p19_s_0__123_comb;
  wire [3:0] p19_s_0__122_comb;
  wire [10:0] p19_s_0__121_comb;
  wire [13:0] p19_s_0__120_comb;
  wire [2:0] p19_s_0__127_comb;
  wire [3:0] p19_s_0__126_comb;
  wire [10:0] p19_s_0__125_comb;
  wire [13:0] p19_s_0__124_comb;
  wire [2:0] p19_s_0__131_comb;
  wire [3:0] p19_s_0__130_comb;
  wire [10:0] p19_s_0__129_comb;
  wire [13:0] p19_s_0__128_comb;
  wire [31:0] p19_temp1__409_comb;
  wire [31:0] p19_value__32_comb;
  wire [31:0] p19_temp2__22_comb;
  wire [31:0] p19_value__47_comb;
  wire [31:0] p19_s_0__18_comb;
  wire [31:0] p19_s_0__19_comb;
  wire [31:0] p19_s_0__20_comb;
  wire [31:0] p19_s_0__21_comb;
  wire [31:0] p19_e__23_comb;
  wire [30:0] p19_add_58872_comb;
  wire [31:0] p19_value__33_comb;
  wire [31:0] p19_a__23_comb;
  wire [31:0] p19_value__48_comb;
  wire [31:0] p19_value__52_comb;
  wire [31:0] p19_value__55_comb;
  wire [31:0] p19_value__58_comb;
  wire [31:0] p19_value__61_comb;
  assign p19_s_1__83_comb = p18_value__21[16:7] ^ p18_value__21[18:9];
  assign p19_s_1__82_comb = p18_value__21[6:0] ^ p18_value__21[8:2] ^ p18_value__21[31:25];
  assign p19_s_1__81_comb = p18_value__21[31:30] ^ p18_value__21[1:0] ^ p18_value__21[24:23];
  assign p19_s_1__80_comb = p18_value__21[29:17] ^ p18_value__21[31:19] ^ p18_value__21[22:10];
  assign p19_S0__147_comb = p18_a__21[1:0] ^ p18_a__21[12:11] ^ p18_a__21[21:20];
  assign p19_S0__146_comb = p18_a__21[31:21] ^ p18_a__21[10:0] ^ p18_a__21[19:9];
  assign p19_S0__145_comb = p18_a__21[20:12] ^ p18_a__21[31:23] ^ p18_a__21[8:0];
  assign p19_S0__144_comb = p18_a__21[11:2] ^ p18_a__21[22:13] ^ p18_a__21[31:22];
  assign p19_and_58906_comb = p18_a__21 & p18_a__20;
  assign p19_s_1__9_comb = {p19_s_1__83_comb, p19_s_1__82_comb, p19_s_1__81_comb, p19_s_1__80_comb};
  assign p19_S0__21_comb = {p19_S0__147_comb, p19_S0__146_comb, p19_S0__145_comb, p19_S0__144_comb};
  assign p19_maj__21_comb = p19_and_58906_comb ^ p18_a__21 & p18_a__19 ^ p18_and_58783;
  assign p19_e__22_comb = p18_a__18 + p18_temp1__412;
  assign p19_value__26_comb = p18_value__6 + p19_s_1__9_comb;
  assign p19_temp2__21_comb = p19_S0__21_comb + p19_maj__21_comb;
  assign p19_value__27_comb = p18_value__25 + p19_value__26_comb;
  assign p19_a__22_comb = p18_temp1__412 + p19_temp2__21_comb;
  assign p19_S1__151_comb = p19_e__22_comb[5:0] ^ p19_e__22_comb[10:5] ^ p19_e__22_comb[24:19];
  assign p19_S1__150_comb = p19_e__22_comb[31:27] ^ p19_e__22_comb[4:0] ^ p19_e__22_comb[18:14];
  assign p19_S1__149_comb = p19_e__22_comb[26:13] ^ p19_e__22_comb[31:18] ^ p19_e__22_comb[13:0];
  assign p19_S1__148_comb = p19_e__22_comb[12:6] ^ p19_e__22_comb[17:11] ^ p19_e__22_comb[31:25];
  assign p19_add_58861_comb = p18_value__21[31:2] + 30'h172c_2a77;
  assign p19_S1__22_comb = {p19_S1__151_comb, p19_S1__150_comb, p19_S1__149_comb, p19_S1__148_comb};
  assign p19_ch__22_comb = p19_e__22_comb & p18_e__21 ^ ~(p19_e__22_comb | ~p18_e__20);
  assign p19_temp1__280_comb = {p19_add_58861_comb, p18_value__21[1:0]};
  assign p19_s_1__91_comb = p19_value__27_comb[16:7] ^ p19_value__27_comb[18:9];
  assign p19_s_1__90_comb = p19_value__27_comb[6:0] ^ p19_value__27_comb[8:2] ^ p19_value__27_comb[31:25];
  assign p19_s_1__89_comb = p19_value__27_comb[31:30] ^ p19_value__27_comb[1:0] ^ p19_value__27_comb[24:23];
  assign p19_s_1__88_comb = p19_value__27_comb[29:17] ^ p19_value__27_comb[31:19] ^ p19_value__27_comb[22:10];
  assign p19_S0__151_comb = p19_a__22_comb[1:0] ^ p19_a__22_comb[12:11] ^ p19_a__22_comb[21:20];
  assign p19_S0__150_comb = p19_a__22_comb[31:21] ^ p19_a__22_comb[10:0] ^ p19_a__22_comb[19:9];
  assign p19_S0__149_comb = p19_a__22_comb[20:12] ^ p19_a__22_comb[31:23] ^ p19_a__22_comb[8:0];
  assign p19_S0__148_comb = p19_a__22_comb[11:2] ^ p19_a__22_comb[22:13] ^ p19_a__22_comb[31:22];
  assign p19_and_58946_comb = p19_a__22_comb & p18_a__21;
  assign p19_s_1__111_comb = p18_value__42[16:7] ^ p18_value__42[18:9];
  assign p19_s_1__110_comb = p18_value__42[6:0] ^ p18_value__42[8:2] ^ p18_value__42[31:25];
  assign p19_s_1__109_comb = p18_value__42[31:30] ^ p18_value__42[1:0] ^ p18_value__42[24:23];
  assign p19_s_1__108_comb = p18_value__42[29:17] ^ p18_value__42[31:19] ^ p18_value__42[22:10];
  assign p19_temp1__407_comb = p18_e__19 + p19_S1__22_comb;
  assign p19_temp1__408_comb = p19_ch__22_comb + p19_temp1__280_comb;
  assign p19_s_1__11_comb = {p19_s_1__91_comb, p19_s_1__90_comb, p19_s_1__89_comb, p19_s_1__88_comb};
  assign p19_S0__22_comb = {p19_S0__151_comb, p19_S0__150_comb, p19_S0__149_comb, p19_S0__148_comb};
  assign p19_maj__22_comb = p19_and_58946_comb ^ p19_a__22_comb & p18_a__20 ^ p19_and_58906_comb;
  assign p19_s_1__16_comb = {p19_s_1__111_comb, p19_s_1__110_comb, p19_s_1__109_comb, p19_s_1__108_comb};
  assign p19_s_0__119_comb = p18_value__9[6:4] ^ p18_value__9[17:15];
  assign p19_s_0__118_comb = p18_value__9[3:0] ^ p18_value__9[14:11] ^ p18_value__9[31:28];
  assign p19_s_0__117_comb = p18_value__9[31:21] ^ p18_value__9[10:0] ^ p18_value__9[27:17];
  assign p19_s_0__116_comb = p18_value__9[20:7] ^ p18_value__9[31:18] ^ p18_value__9[16:3];
  assign p19_s_0__123_comb = p18_value__12[6:4] ^ p18_value__12[17:15];
  assign p19_s_0__122_comb = p18_value__12[3:0] ^ p18_value__12[14:11] ^ p18_value__12[31:28];
  assign p19_s_0__121_comb = p18_value__12[31:21] ^ p18_value__12[10:0] ^ p18_value__12[27:17];
  assign p19_s_0__120_comb = p18_value__12[20:7] ^ p18_value__12[31:18] ^ p18_value__12[16:3];
  assign p19_s_0__127_comb = p18_value__15[6:4] ^ p18_value__15[17:15];
  assign p19_s_0__126_comb = p18_value__15[3:0] ^ p18_value__15[14:11] ^ p18_value__15[31:28];
  assign p19_s_0__125_comb = p18_value__15[31:21] ^ p18_value__15[10:0] ^ p18_value__15[27:17];
  assign p19_s_0__124_comb = p18_value__15[20:7] ^ p18_value__15[31:18] ^ p18_value__15[16:3];
  assign p19_s_0__131_comb = p18_value__18[6:4] ^ p18_value__18[17:15];
  assign p19_s_0__130_comb = p18_value__18[3:0] ^ p18_value__18[14:11] ^ p18_value__18[31:28];
  assign p19_s_0__129_comb = p18_value__18[31:21] ^ p18_value__18[10:0] ^ p18_value__18[27:17];
  assign p19_s_0__128_comb = p18_value__18[20:7] ^ p18_value__18[31:18] ^ p18_value__18[16:3];
  assign p19_temp1__409_comb = p19_temp1__407_comb + p19_temp1__408_comb;
  assign p19_value__32_comb = p18_value__12 + p19_s_1__11_comb;
  assign p19_temp2__22_comb = p19_S0__22_comb + p19_maj__22_comb;
  assign p19_value__47_comb = p19_value__27_comb + p19_s_1__16_comb;
  assign p19_s_0__18_comb = {p19_s_0__119_comb, p19_s_0__118_comb, p19_s_0__117_comb, p19_s_0__116_comb};
  assign p19_s_0__19_comb = {p19_s_0__123_comb, p19_s_0__122_comb, p19_s_0__121_comb, p19_s_0__120_comb};
  assign p19_s_0__20_comb = {p19_s_0__127_comb, p19_s_0__126_comb, p19_s_0__125_comb, p19_s_0__124_comb};
  assign p19_s_0__21_comb = {p19_s_0__131_comb, p19_s_0__130_comb, p19_s_0__129_comb, p19_s_0__128_comb};
  assign p19_e__23_comb = p18_a__19 + p19_temp1__409_comb;
  assign p19_add_58872_comb = p18_value__24[31:1] + 31'h3b7c_c46d;
  assign p19_value__33_comb = p18_value__31 + p19_value__32_comb;
  assign p19_a__23_comb = p19_temp1__409_comb + p19_temp2__22_comb;
  assign p19_value__48_comb = p18_value__46 + p19_value__47_comb;
  assign p19_value__52_comb = p18_value__6 + p19_s_0__18_comb;
  assign p19_value__55_comb = p18_value__9 + p19_s_0__19_comb;
  assign p19_value__58_comb = p18_value__12 + p19_s_0__20_comb;
  assign p19_value__61_comb = p18_value__15 + p19_s_0__21_comb;

  // Registers for pipe stage 19:
  reg [31:0] p19_e__20;
  reg [31:0] p19_e__21;
  reg [31:0] p19_value__18;
  reg [31:0] p19_e__22;
  reg [31:0] p19_value__21;
  reg [31:0] p19_e__23;
  reg [31:0] p19_value__24;
  reg [30:0] p19_add_58872;
  reg [31:0] p19_a__20;
  reg [31:0] p19_value__27;
  reg [31:0] p19_a__21;
  reg [31:0] p19_value__30;
  reg [31:0] p19_a__22;
  reg [31:0] p19_value__33;
  reg [31:0] p19_and_58946;
  reg [31:0] p19_a__23;
  reg [31:0] p19_value__36;
  reg [31:0] p19_value__37;
  reg [31:0] p19_value__42;
  reg [31:0] p19_value__43;
  reg [31:0] p19_value__48;
  reg [31:0] p19_value__49;
  reg [31:0] p19_value__52;
  reg [31:0] p19_value__55;
  reg [31:0] p19_value__58;
  reg [31:0] p19_value__61;
  always_ff @ (posedge clk) begin
    p19_e__20 <= p18_e__20;
    p19_e__21 <= p18_e__21;
    p19_value__18 <= p18_value__18;
    p19_e__22 <= p19_e__22_comb;
    p19_value__21 <= p18_value__21;
    p19_e__23 <= p19_e__23_comb;
    p19_value__24 <= p18_value__24;
    p19_add_58872 <= p19_add_58872_comb;
    p19_a__20 <= p18_a__20;
    p19_value__27 <= p19_value__27_comb;
    p19_a__21 <= p18_a__21;
    p19_value__30 <= p18_value__30;
    p19_a__22 <= p19_a__22_comb;
    p19_value__33 <= p19_value__33_comb;
    p19_and_58946 <= p19_and_58946_comb;
    p19_a__23 <= p19_a__23_comb;
    p19_value__36 <= p18_value__36;
    p19_value__37 <= p18_value__37;
    p19_value__42 <= p18_value__42;
    p19_value__43 <= p18_value__43;
    p19_value__48 <= p19_value__48_comb;
    p19_value__49 <= p18_value__49;
    p19_value__52 <= p19_value__52_comb;
    p19_value__55 <= p19_value__55_comb;
    p19_value__58 <= p19_value__58_comb;
    p19_value__61 <= p19_value__61_comb;
  end

  // ===== Pipe stage 20:
  wire [5:0] p20_S1__155_comb;
  wire [4:0] p20_S1__154_comb;
  wire [13:0] p20_S1__153_comb;
  wire [6:0] p20_S1__152_comb;
  wire [9:0] p20_s_1__99_comb;
  wire [6:0] p20_s_1__98_comb;
  wire [1:0] p20_s_1__97_comb;
  wire [12:0] p20_s_1__96_comb;
  wire [9:0] p20_s_1__119_comb;
  wire [6:0] p20_s_1__118_comb;
  wire [1:0] p20_s_1__117_comb;
  wire [12:0] p20_s_1__116_comb;
  wire [31:0] p20_S1__23_comb;
  wire [31:0] p20_ch__23_comb;
  wire [31:0] p20_temp1__281_comb;
  wire [31:0] p20_s_1__13_comb;
  wire [31:0] p20_s_1__18_comb;
  wire [31:0] p20_temp1__404_comb;
  wire [31:0] p20_temp1__405_comb;
  wire [31:0] p20_value__38_comb;
  wire [31:0] p20_value__53_comb;
  wire [31:0] p20_temp1__406_comb;
  wire [31:0] p20_value__39_comb;
  wire [31:0] p20_value__54_comb;
  wire [31:0] p20_e__24_comb;
  wire [1:0] p20_S0__155_comb;
  wire [10:0] p20_S0__154_comb;
  wire [8:0] p20_S0__153_comb;
  wire [9:0] p20_S0__152_comb;
  wire [31:0] p20_and_59161_comb;
  wire [9:0] p20_s_1__107_comb;
  wire [6:0] p20_s_1__106_comb;
  wire [1:0] p20_s_1__105_comb;
  wire [12:0] p20_s_1__104_comb;
  wire [9:0] p20_s_1__127_comb;
  wire [6:0] p20_s_1__126_comb;
  wire [1:0] p20_s_1__125_comb;
  wire [12:0] p20_s_1__124_comb;
  wire [5:0] p20_S1__159_comb;
  wire [4:0] p20_S1__158_comb;
  wire [13:0] p20_S1__157_comb;
  wire [6:0] p20_S1__156_comb;
  wire [30:0] p20_add_59138_comb;
  wire [31:0] p20_S0__23_comb;
  wire [31:0] p20_maj__23_comb;
  wire [31:0] p20_s_1__15_comb;
  wire [31:0] p20_s_1__20_comb;
  wire [2:0] p20_s_0__135_comb;
  wire [3:0] p20_s_0__134_comb;
  wire [10:0] p20_s_0__133_comb;
  wire [13:0] p20_s_0__132_comb;
  wire [2:0] p20_s_0__139_comb;
  wire [3:0] p20_s_0__138_comb;
  wire [10:0] p20_s_0__137_comb;
  wire [13:0] p20_s_0__136_comb;
  wire [2:0] p20_s_0__143_comb;
  wire [3:0] p20_s_0__142_comb;
  wire [10:0] p20_s_0__141_comb;
  wire [13:0] p20_s_0__140_comb;
  wire [2:0] p20_s_0__147_comb;
  wire [3:0] p20_s_0__146_comb;
  wire [10:0] p20_s_0__145_comb;
  wire [13:0] p20_s_0__144_comb;
  wire [31:0] p20_S1__24_comb;
  wire [31:0] p20_ch__24_comb;
  wire [31:0] p20_temp1__282_comb;
  wire [31:0] p20_temp2__23_comb;
  wire [31:0] p20_value__44_comb;
  wire [31:0] p20_value__59_comb;
  wire [31:0] p20_s_0__22_comb;
  wire [31:0] p20_s_0__23_comb;
  wire [31:0] p20_s_0__24_comb;
  wire [31:0] p20_s_0__25_comb;
  wire [31:0] p20_temp1__401_comb;
  wire [31:0] p20_temp1__402_comb;
  wire [31:0] p20_a__24_comb;
  wire [31:0] p20_value__45_comb;
  wire [31:0] p20_value__60_comb;
  wire [31:0] p20_value__64_comb;
  wire [31:0] p20_value__67_comb;
  wire [31:0] p20_value__70_comb;
  wire [31:0] p20_value__73_comb;
  assign p20_S1__155_comb = p19_e__23[5:0] ^ p19_e__23[10:5] ^ p19_e__23[24:19];
  assign p20_S1__154_comb = p19_e__23[31:27] ^ p19_e__23[4:0] ^ p19_e__23[18:14];
  assign p20_S1__153_comb = p19_e__23[26:13] ^ p19_e__23[31:18] ^ p19_e__23[13:0];
  assign p20_S1__152_comb = p19_e__23[12:6] ^ p19_e__23[17:11] ^ p19_e__23[31:25];
  assign p20_s_1__99_comb = p19_value__33[16:7] ^ p19_value__33[18:9];
  assign p20_s_1__98_comb = p19_value__33[6:0] ^ p19_value__33[8:2] ^ p19_value__33[31:25];
  assign p20_s_1__97_comb = p19_value__33[31:30] ^ p19_value__33[1:0] ^ p19_value__33[24:23];
  assign p20_s_1__96_comb = p19_value__33[29:17] ^ p19_value__33[31:19] ^ p19_value__33[22:10];
  assign p20_s_1__119_comb = p19_value__48[16:7] ^ p19_value__48[18:9];
  assign p20_s_1__118_comb = p19_value__48[6:0] ^ p19_value__48[8:2] ^ p19_value__48[31:25];
  assign p20_s_1__117_comb = p19_value__48[31:30] ^ p19_value__48[1:0] ^ p19_value__48[24:23];
  assign p20_s_1__116_comb = p19_value__48[29:17] ^ p19_value__48[31:19] ^ p19_value__48[22:10];
  assign p20_S1__23_comb = {p20_S1__155_comb, p20_S1__154_comb, p20_S1__153_comb, p20_S1__152_comb};
  assign p20_ch__23_comb = p19_e__23 & p19_e__22 ^ ~(p19_e__23 | ~p19_e__21);
  assign p20_temp1__281_comb = {p19_add_58872, p19_value__24[0]};
  assign p20_s_1__13_comb = {p20_s_1__99_comb, p20_s_1__98_comb, p20_s_1__97_comb, p20_s_1__96_comb};
  assign p20_s_1__18_comb = {p20_s_1__119_comb, p20_s_1__118_comb, p20_s_1__117_comb, p20_s_1__116_comb};
  assign p20_temp1__404_comb = p19_e__20 + p20_S1__23_comb;
  assign p20_temp1__405_comb = p20_ch__23_comb + p20_temp1__281_comb;
  assign p20_value__38_comb = p19_value__18 + p20_s_1__13_comb;
  assign p20_value__53_comb = p19_value__33 + p20_s_1__18_comb;
  assign p20_temp1__406_comb = p20_temp1__404_comb + p20_temp1__405_comb;
  assign p20_value__39_comb = p19_value__37 + p20_value__38_comb;
  assign p20_value__54_comb = p19_value__52 + p20_value__53_comb;
  assign p20_e__24_comb = p19_a__20 + p20_temp1__406_comb;
  assign p20_S0__155_comb = p19_a__23[1:0] ^ p19_a__23[12:11] ^ p19_a__23[21:20];
  assign p20_S0__154_comb = p19_a__23[31:21] ^ p19_a__23[10:0] ^ p19_a__23[19:9];
  assign p20_S0__153_comb = p19_a__23[20:12] ^ p19_a__23[31:23] ^ p19_a__23[8:0];
  assign p20_S0__152_comb = p19_a__23[11:2] ^ p19_a__23[22:13] ^ p19_a__23[31:22];
  assign p20_and_59161_comb = p19_a__23 & p19_a__22;
  assign p20_s_1__107_comb = p20_value__39_comb[16:7] ^ p20_value__39_comb[18:9];
  assign p20_s_1__106_comb = p20_value__39_comb[6:0] ^ p20_value__39_comb[8:2] ^ p20_value__39_comb[31:25];
  assign p20_s_1__105_comb = p20_value__39_comb[31:30] ^ p20_value__39_comb[1:0] ^ p20_value__39_comb[24:23];
  assign p20_s_1__104_comb = p20_value__39_comb[29:17] ^ p20_value__39_comb[31:19] ^ p20_value__39_comb[22:10];
  assign p20_s_1__127_comb = p20_value__54_comb[16:7] ^ p20_value__54_comb[18:9];
  assign p20_s_1__126_comb = p20_value__54_comb[6:0] ^ p20_value__54_comb[8:2] ^ p20_value__54_comb[31:25];
  assign p20_s_1__125_comb = p20_value__54_comb[31:30] ^ p20_value__54_comb[1:0] ^ p20_value__54_comb[24:23];
  assign p20_s_1__124_comb = p20_value__54_comb[29:17] ^ p20_value__54_comb[31:19] ^ p20_value__54_comb[22:10];
  assign p20_S1__159_comb = p20_e__24_comb[5:0] ^ p20_e__24_comb[10:5] ^ p20_e__24_comb[24:19];
  assign p20_S1__158_comb = p20_e__24_comb[31:27] ^ p20_e__24_comb[4:0] ^ p20_e__24_comb[18:14];
  assign p20_S1__157_comb = p20_e__24_comb[26:13] ^ p20_e__24_comb[31:18] ^ p20_e__24_comb[13:0];
  assign p20_S1__156_comb = p20_e__24_comb[12:6] ^ p20_e__24_comb[17:11] ^ p20_e__24_comb[31:25];
  assign p20_add_59138_comb = p19_value__27[31:1] + 31'h4c1f_28a9;
  assign p20_S0__23_comb = {p20_S0__155_comb, p20_S0__154_comb, p20_S0__153_comb, p20_S0__152_comb};
  assign p20_maj__23_comb = p20_and_59161_comb ^ p19_a__23 & p19_a__21 ^ p19_and_58946;
  assign p20_s_1__15_comb = {p20_s_1__107_comb, p20_s_1__106_comb, p20_s_1__105_comb, p20_s_1__104_comb};
  assign p20_s_1__20_comb = {p20_s_1__127_comb, p20_s_1__126_comb, p20_s_1__125_comb, p20_s_1__124_comb};
  assign p20_s_0__135_comb = p19_value__21[6:4] ^ p19_value__21[17:15];
  assign p20_s_0__134_comb = p19_value__21[3:0] ^ p19_value__21[14:11] ^ p19_value__21[31:28];
  assign p20_s_0__133_comb = p19_value__21[31:21] ^ p19_value__21[10:0] ^ p19_value__21[27:17];
  assign p20_s_0__132_comb = p19_value__21[20:7] ^ p19_value__21[31:18] ^ p19_value__21[16:3];
  assign p20_s_0__139_comb = p19_value__24[6:4] ^ p19_value__24[17:15];
  assign p20_s_0__138_comb = p19_value__24[3:0] ^ p19_value__24[14:11] ^ p19_value__24[31:28];
  assign p20_s_0__137_comb = p19_value__24[31:21] ^ p19_value__24[10:0] ^ p19_value__24[27:17];
  assign p20_s_0__136_comb = p19_value__24[20:7] ^ p19_value__24[31:18] ^ p19_value__24[16:3];
  assign p20_s_0__143_comb = p19_value__27[6:4] ^ p19_value__27[17:15];
  assign p20_s_0__142_comb = p19_value__27[3:0] ^ p19_value__27[14:11] ^ p19_value__27[31:28];
  assign p20_s_0__141_comb = p19_value__27[31:21] ^ p19_value__27[10:0] ^ p19_value__27[27:17];
  assign p20_s_0__140_comb = p19_value__27[20:7] ^ p19_value__27[31:18] ^ p19_value__27[16:3];
  assign p20_s_0__147_comb = p19_value__30[6:4] ^ p19_value__30[17:15];
  assign p20_s_0__146_comb = p19_value__30[3:0] ^ p19_value__30[14:11] ^ p19_value__30[31:28];
  assign p20_s_0__145_comb = p19_value__30[31:21] ^ p19_value__30[10:0] ^ p19_value__30[27:17];
  assign p20_s_0__144_comb = p19_value__30[20:7] ^ p19_value__30[31:18] ^ p19_value__30[16:3];
  assign p20_S1__24_comb = {p20_S1__159_comb, p20_S1__158_comb, p20_S1__157_comb, p20_S1__156_comb};
  assign p20_ch__24_comb = p20_e__24_comb & p19_e__23 ^ ~(p20_e__24_comb | ~p19_e__22);
  assign p20_temp1__282_comb = {p20_add_59138_comb, p19_value__27[0]};
  assign p20_temp2__23_comb = p20_S0__23_comb + p20_maj__23_comb;
  assign p20_value__44_comb = p19_value__24 + p20_s_1__15_comb;
  assign p20_value__59_comb = p20_value__39_comb + p20_s_1__20_comb;
  assign p20_s_0__22_comb = {p20_s_0__135_comb, p20_s_0__134_comb, p20_s_0__133_comb, p20_s_0__132_comb};
  assign p20_s_0__23_comb = {p20_s_0__139_comb, p20_s_0__138_comb, p20_s_0__137_comb, p20_s_0__136_comb};
  assign p20_s_0__24_comb = {p20_s_0__143_comb, p20_s_0__142_comb, p20_s_0__141_comb, p20_s_0__140_comb};
  assign p20_s_0__25_comb = {p20_s_0__147_comb, p20_s_0__146_comb, p20_s_0__145_comb, p20_s_0__144_comb};
  assign p20_temp1__401_comb = p19_e__21 + p20_S1__24_comb;
  assign p20_temp1__402_comb = p20_ch__24_comb + p20_temp1__282_comb;
  assign p20_a__24_comb = p20_temp1__406_comb + p20_temp2__23_comb;
  assign p20_value__45_comb = p19_value__43 + p20_value__44_comb;
  assign p20_value__60_comb = p19_value__58 + p20_value__59_comb;
  assign p20_value__64_comb = p19_value__18 + p20_s_0__22_comb;
  assign p20_value__67_comb = p19_value__21 + p20_s_0__23_comb;
  assign p20_value__70_comb = p19_value__24 + p20_s_0__24_comb;
  assign p20_value__73_comb = p19_value__27 + p20_s_0__25_comb;

  // Registers for pipe stage 20:
  reg [31:0] p20_e__22;
  reg [31:0] p20_e__23;
  reg [31:0] p20_e__24;
  reg [31:0] p20_temp1__401;
  reg [31:0] p20_temp1__402;
  reg [31:0] p20_a__21;
  reg [31:0] p20_value__30;
  reg [31:0] p20_a__22;
  reg [31:0] p20_value__33;
  reg [31:0] p20_a__23;
  reg [31:0] p20_and_59161;
  reg [31:0] p20_value__36;
  reg [31:0] p20_a__24;
  reg [31:0] p20_value__39;
  reg [31:0] p20_value__42;
  reg [31:0] p20_value__45;
  reg [31:0] p20_value__48;
  reg [31:0] p20_value__49;
  reg [31:0] p20_value__54;
  reg [31:0] p20_value__55;
  reg [31:0] p20_value__60;
  reg [31:0] p20_value__61;
  reg [31:0] p20_value__64;
  reg [31:0] p20_value__67;
  reg [31:0] p20_value__70;
  reg [31:0] p20_value__73;
  always_ff @ (posedge clk) begin
    p20_e__22 <= p19_e__22;
    p20_e__23 <= p19_e__23;
    p20_e__24 <= p20_e__24_comb;
    p20_temp1__401 <= p20_temp1__401_comb;
    p20_temp1__402 <= p20_temp1__402_comb;
    p20_a__21 <= p19_a__21;
    p20_value__30 <= p19_value__30;
    p20_a__22 <= p19_a__22;
    p20_value__33 <= p19_value__33;
    p20_a__23 <= p19_a__23;
    p20_and_59161 <= p20_and_59161_comb;
    p20_value__36 <= p19_value__36;
    p20_a__24 <= p20_a__24_comb;
    p20_value__39 <= p20_value__39_comb;
    p20_value__42 <= p19_value__42;
    p20_value__45 <= p20_value__45_comb;
    p20_value__48 <= p19_value__48;
    p20_value__49 <= p19_value__49;
    p20_value__54 <= p20_value__54_comb;
    p20_value__55 <= p19_value__55;
    p20_value__60 <= p20_value__60_comb;
    p20_value__61 <= p19_value__61;
    p20_value__64 <= p20_value__64_comb;
    p20_value__67 <= p20_value__67_comb;
    p20_value__70 <= p20_value__70_comb;
    p20_value__73 <= p20_value__73_comb;
  end

  // ===== Pipe stage 21:
  wire [9:0] p21_s_1__115_comb;
  wire [6:0] p21_s_1__114_comb;
  wire [1:0] p21_s_1__113_comb;
  wire [12:0] p21_s_1__112_comb;
  wire [9:0] p21_s_1__135_comb;
  wire [6:0] p21_s_1__134_comb;
  wire [1:0] p21_s_1__133_comb;
  wire [12:0] p21_s_1__132_comb;
  wire [31:0] p21_s_1__17_comb;
  wire [31:0] p21_s_1__22_comb;
  wire [31:0] p21_temp1__403_comb;
  wire [31:0] p21_value__50_comb;
  wire [31:0] p21_value__65_comb;
  wire [31:0] p21_e__25_comb;
  wire [31:0] p21_value__51_comb;
  wire [31:0] p21_value__66_comb;
  wire [5:0] p21_S1__163_comb;
  wire [4:0] p21_S1__162_comb;
  wire [13:0] p21_S1__161_comb;
  wire [6:0] p21_S1__160_comb;
  wire [1:0] p21_S0__159_comb;
  wire [10:0] p21_S0__158_comb;
  wire [8:0] p21_S0__157_comb;
  wire [9:0] p21_S0__156_comb;
  wire [31:0] p21_and_59402_comb;
  wire [9:0] p21_s_1__123_comb;
  wire [6:0] p21_s_1__122_comb;
  wire [1:0] p21_s_1__121_comb;
  wire [12:0] p21_s_1__120_comb;
  wire [9:0] p21_s_1__143_comb;
  wire [6:0] p21_s_1__142_comb;
  wire [1:0] p21_s_1__141_comb;
  wire [12:0] p21_s_1__140_comb;
  wire [31:0] p21_S1__25_comb;
  wire [31:0] p21_S0__24_comb;
  wire [31:0] p21_maj__24_comb;
  wire [31:0] p21_s_1__19_comb;
  wire [31:0] p21_s_1__24_comb;
  wire [2:0] p21_s_0__151_comb;
  wire [3:0] p21_s_0__150_comb;
  wire [10:0] p21_s_0__149_comb;
  wire [13:0] p21_s_0__148_comb;
  wire [31:0] p21_temp1__101_comb;
  wire [31:0] p21_ch__25_comb;
  wire [31:0] p21_temp2__24_comb;
  wire [31:0] p21_value__56_comb;
  wire [31:0] p21_value__71_comb;
  wire [31:0] p21_s_0__26_comb;
  wire [31:0] p21_temp1__102_comb;
  wire [31:0] p21_temp1__283_comb;
  wire [31:0] p21_a__25_comb;
  wire [31:0] p21_value__57_comb;
  wire [31:0] p21_value__72_comb;
  wire [31:0] p21_value__76_comb;
  assign p21_s_1__115_comb = p20_value__45[16:7] ^ p20_value__45[18:9];
  assign p21_s_1__114_comb = p20_value__45[6:0] ^ p20_value__45[8:2] ^ p20_value__45[31:25];
  assign p21_s_1__113_comb = p20_value__45[31:30] ^ p20_value__45[1:0] ^ p20_value__45[24:23];
  assign p21_s_1__112_comb = p20_value__45[29:17] ^ p20_value__45[31:19] ^ p20_value__45[22:10];
  assign p21_s_1__135_comb = p20_value__60[16:7] ^ p20_value__60[18:9];
  assign p21_s_1__134_comb = p20_value__60[6:0] ^ p20_value__60[8:2] ^ p20_value__60[31:25];
  assign p21_s_1__133_comb = p20_value__60[31:30] ^ p20_value__60[1:0] ^ p20_value__60[24:23];
  assign p21_s_1__132_comb = p20_value__60[29:17] ^ p20_value__60[31:19] ^ p20_value__60[22:10];
  assign p21_s_1__17_comb = {p21_s_1__115_comb, p21_s_1__114_comb, p21_s_1__113_comb, p21_s_1__112_comb};
  assign p21_s_1__22_comb = {p21_s_1__135_comb, p21_s_1__134_comb, p21_s_1__133_comb, p21_s_1__132_comb};
  assign p21_temp1__403_comb = p20_temp1__401 + p20_temp1__402;
  assign p21_value__50_comb = p20_value__30 + p21_s_1__17_comb;
  assign p21_value__65_comb = p20_value__45 + p21_s_1__22_comb;
  assign p21_e__25_comb = p20_a__21 + p21_temp1__403_comb;
  assign p21_value__51_comb = p20_value__49 + p21_value__50_comb;
  assign p21_value__66_comb = p20_value__64 + p21_value__65_comb;
  assign p21_S1__163_comb = p21_e__25_comb[5:0] ^ p21_e__25_comb[10:5] ^ p21_e__25_comb[24:19];
  assign p21_S1__162_comb = p21_e__25_comb[31:27] ^ p21_e__25_comb[4:0] ^ p21_e__25_comb[18:14];
  assign p21_S1__161_comb = p21_e__25_comb[26:13] ^ p21_e__25_comb[31:18] ^ p21_e__25_comb[13:0];
  assign p21_S1__160_comb = p21_e__25_comb[12:6] ^ p21_e__25_comb[17:11] ^ p21_e__25_comb[31:25];
  assign p21_S0__159_comb = p20_a__24[1:0] ^ p20_a__24[12:11] ^ p20_a__24[21:20];
  assign p21_S0__158_comb = p20_a__24[31:21] ^ p20_a__24[10:0] ^ p20_a__24[19:9];
  assign p21_S0__157_comb = p20_a__24[20:12] ^ p20_a__24[31:23] ^ p20_a__24[8:0];
  assign p21_S0__156_comb = p20_a__24[11:2] ^ p20_a__24[22:13] ^ p20_a__24[31:22];
  assign p21_and_59402_comb = p20_a__24 & p20_a__23;
  assign p21_s_1__123_comb = p21_value__51_comb[16:7] ^ p21_value__51_comb[18:9];
  assign p21_s_1__122_comb = p21_value__51_comb[6:0] ^ p21_value__51_comb[8:2] ^ p21_value__51_comb[31:25];
  assign p21_s_1__121_comb = p21_value__51_comb[31:30] ^ p21_value__51_comb[1:0] ^ p21_value__51_comb[24:23];
  assign p21_s_1__120_comb = p21_value__51_comb[29:17] ^ p21_value__51_comb[31:19] ^ p21_value__51_comb[22:10];
  assign p21_s_1__143_comb = p21_value__66_comb[16:7] ^ p21_value__66_comb[18:9];
  assign p21_s_1__142_comb = p21_value__66_comb[6:0] ^ p21_value__66_comb[8:2] ^ p21_value__66_comb[31:25];
  assign p21_s_1__141_comb = p21_value__66_comb[31:30] ^ p21_value__66_comb[1:0] ^ p21_value__66_comb[24:23];
  assign p21_s_1__140_comb = p21_value__66_comb[29:17] ^ p21_value__66_comb[31:19] ^ p21_value__66_comb[22:10];
  assign p21_S1__25_comb = {p21_S1__163_comb, p21_S1__162_comb, p21_S1__161_comb, p21_S1__160_comb};
  assign p21_S0__24_comb = {p21_S0__159_comb, p21_S0__158_comb, p21_S0__157_comb, p21_S0__156_comb};
  assign p21_maj__24_comb = p21_and_59402_comb ^ p20_a__24 & p20_a__22 ^ p20_and_59161;
  assign p21_s_1__19_comb = {p21_s_1__123_comb, p21_s_1__122_comb, p21_s_1__121_comb, p21_s_1__120_comb};
  assign p21_s_1__24_comb = {p21_s_1__143_comb, p21_s_1__142_comb, p21_s_1__141_comb, p21_s_1__140_comb};
  assign p21_s_0__151_comb = p20_value__33[6:4] ^ p20_value__33[17:15];
  assign p21_s_0__150_comb = p20_value__33[3:0] ^ p20_value__33[14:11] ^ p20_value__33[31:28];
  assign p21_s_0__149_comb = p20_value__33[31:21] ^ p20_value__33[10:0] ^ p20_value__33[27:17];
  assign p21_s_0__148_comb = p20_value__33[20:7] ^ p20_value__33[31:18] ^ p20_value__33[16:3];
  assign p21_temp1__101_comb = p20_e__22 + p21_S1__25_comb;
  assign p21_ch__25_comb = p21_e__25_comb & p20_e__24 ^ ~(p21_e__25_comb | ~p20_e__23);
  assign p21_temp2__24_comb = p21_S0__24_comb + p21_maj__24_comb;
  assign p21_value__56_comb = p20_value__36 + p21_s_1__19_comb;
  assign p21_value__71_comb = p21_value__51_comb + p21_s_1__24_comb;
  assign p21_s_0__26_comb = {p21_s_0__151_comb, p21_s_0__150_comb, p21_s_0__149_comb, p21_s_0__148_comb};
  assign p21_temp1__102_comb = p21_temp1__101_comb + p21_ch__25_comb;
  assign p21_temp1__283_comb = p20_value__30 + 32'ha831_c66d;
  assign p21_a__25_comb = p21_temp1__403_comb + p21_temp2__24_comb;
  assign p21_value__57_comb = p20_value__55 + p21_value__56_comb;
  assign p21_value__72_comb = p20_value__70 + p21_value__71_comb;
  assign p21_value__76_comb = p20_value__30 + p21_s_0__26_comb;

  // Registers for pipe stage 21:
  reg [31:0] p21_e__23;
  reg [31:0] p21_e__24;
  reg [31:0] p21_e__25;
  reg [31:0] p21_temp1__102;
  reg [31:0] p21_temp1__283;
  reg [31:0] p21_a__22;
  reg [31:0] p21_value__33;
  reg [31:0] p21_a__23;
  reg [31:0] p21_value__36;
  reg [31:0] p21_a__24;
  reg [31:0] p21_and_59402;
  reg [31:0] p21_value__39;
  reg [31:0] p21_a__25;
  reg [31:0] p21_value__42;
  reg [31:0] p21_value__45;
  reg [31:0] p21_value__48;
  reg [31:0] p21_value__51;
  reg [31:0] p21_value__54;
  reg [31:0] p21_value__57;
  reg [31:0] p21_value__60;
  reg [31:0] p21_value__61;
  reg [31:0] p21_value__66;
  reg [31:0] p21_value__67;
  reg [31:0] p21_value__72;
  reg [31:0] p21_value__73;
  reg [31:0] p21_value__76;
  always_ff @ (posedge clk) begin
    p21_e__23 <= p20_e__23;
    p21_e__24 <= p20_e__24;
    p21_e__25 <= p21_e__25_comb;
    p21_temp1__102 <= p21_temp1__102_comb;
    p21_temp1__283 <= p21_temp1__283_comb;
    p21_a__22 <= p20_a__22;
    p21_value__33 <= p20_value__33;
    p21_a__23 <= p20_a__23;
    p21_value__36 <= p20_value__36;
    p21_a__24 <= p20_a__24;
    p21_and_59402 <= p21_and_59402_comb;
    p21_value__39 <= p20_value__39;
    p21_a__25 <= p21_a__25_comb;
    p21_value__42 <= p20_value__42;
    p21_value__45 <= p20_value__45;
    p21_value__48 <= p20_value__48;
    p21_value__51 <= p21_value__51_comb;
    p21_value__54 <= p20_value__54;
    p21_value__57 <= p21_value__57_comb;
    p21_value__60 <= p20_value__60;
    p21_value__61 <= p20_value__61;
    p21_value__66 <= p21_value__66_comb;
    p21_value__67 <= p20_value__67;
    p21_value__72 <= p21_value__72_comb;
    p21_value__73 <= p20_value__73;
    p21_value__76 <= p21_value__76_comb;
  end

  // ===== Pipe stage 22:
  wire [31:0] p22_temp1__104_comb;
  wire [31:0] p22_e__26_comb;
  wire [5:0] p22_S1__167_comb;
  wire [4:0] p22_S1__166_comb;
  wire [13:0] p22_S1__165_comb;
  wire [6:0] p22_S1__164_comb;
  wire [28:0] p22_add_59572_comb;
  wire [1:0] p22_S0__163_comb;
  wire [10:0] p22_S0__162_comb;
  wire [8:0] p22_S0__161_comb;
  wire [9:0] p22_S0__160_comb;
  wire [31:0] p22_and_59596_comb;
  wire [9:0] p22_s_1__151_comb;
  wire [6:0] p22_s_1__150_comb;
  wire [1:0] p22_s_1__149_comb;
  wire [12:0] p22_s_1__148_comb;
  wire [31:0] p22_S1__26_comb;
  wire [31:0] p22_ch__26_comb;
  wire [31:0] p22_temp1__284_comb;
  wire [31:0] p22_S0__25_comb;
  wire [31:0] p22_maj__25_comb;
  wire [31:0] p22_s_1__26_comb;
  wire [2:0] p22_s_0__155_comb;
  wire [3:0] p22_s_0__154_comb;
  wire [10:0] p22_s_0__153_comb;
  wire [13:0] p22_s_0__152_comb;
  wire [31:0] p22_temp1__398_comb;
  wire [31:0] p22_temp1__399_comb;
  wire [31:0] p22_temp2__25_comb;
  wire [31:0] p22_value__77_comb;
  wire [31:0] p22_s_0__27_comb;
  wire [31:0] p22_temp1__400_comb;
  wire [31:0] p22_a__26_comb;
  wire [31:0] p22_value__78_comb;
  wire [31:0] p22_value__79_comb;
  assign p22_temp1__104_comb = p21_temp1__102 + p21_temp1__283;
  assign p22_e__26_comb = p21_a__22 + p22_temp1__104_comb;
  assign p22_S1__167_comb = p22_e__26_comb[5:0] ^ p22_e__26_comb[10:5] ^ p22_e__26_comb[24:19];
  assign p22_S1__166_comb = p22_e__26_comb[31:27] ^ p22_e__26_comb[4:0] ^ p22_e__26_comb[18:14];
  assign p22_S1__165_comb = p22_e__26_comb[26:13] ^ p22_e__26_comb[31:18] ^ p22_e__26_comb[13:0];
  assign p22_S1__164_comb = p22_e__26_comb[12:6] ^ p22_e__26_comb[17:11] ^ p22_e__26_comb[31:25];
  assign p22_add_59572_comb = p21_value__33[31:3] + 29'h1600_64f9;
  assign p22_S0__163_comb = p21_a__25[1:0] ^ p21_a__25[12:11] ^ p21_a__25[21:20];
  assign p22_S0__162_comb = p21_a__25[31:21] ^ p21_a__25[10:0] ^ p21_a__25[19:9];
  assign p22_S0__161_comb = p21_a__25[20:12] ^ p21_a__25[31:23] ^ p21_a__25[8:0];
  assign p22_S0__160_comb = p21_a__25[11:2] ^ p21_a__25[22:13] ^ p21_a__25[31:22];
  assign p22_and_59596_comb = p21_a__25 & p21_a__24;
  assign p22_s_1__151_comb = p21_value__72[16:7] ^ p21_value__72[18:9];
  assign p22_s_1__150_comb = p21_value__72[6:0] ^ p21_value__72[8:2] ^ p21_value__72[31:25];
  assign p22_s_1__149_comb = p21_value__72[31:30] ^ p21_value__72[1:0] ^ p21_value__72[24:23];
  assign p22_s_1__148_comb = p21_value__72[29:17] ^ p21_value__72[31:19] ^ p21_value__72[22:10];
  assign p22_S1__26_comb = {p22_S1__167_comb, p22_S1__166_comb, p22_S1__165_comb, p22_S1__164_comb};
  assign p22_ch__26_comb = p22_e__26_comb & p21_e__25 ^ ~(p22_e__26_comb | ~p21_e__24);
  assign p22_temp1__284_comb = {p22_add_59572_comb, p21_value__33[2:0]};
  assign p22_S0__25_comb = {p22_S0__163_comb, p22_S0__162_comb, p22_S0__161_comb, p22_S0__160_comb};
  assign p22_maj__25_comb = p22_and_59596_comb ^ p21_a__25 & p21_a__23 ^ p21_and_59402;
  assign p22_s_1__26_comb = {p22_s_1__151_comb, p22_s_1__150_comb, p22_s_1__149_comb, p22_s_1__148_comb};
  assign p22_s_0__155_comb = p21_value__36[6:4] ^ p21_value__36[17:15];
  assign p22_s_0__154_comb = p21_value__36[3:0] ^ p21_value__36[14:11] ^ p21_value__36[31:28];
  assign p22_s_0__153_comb = p21_value__36[31:21] ^ p21_value__36[10:0] ^ p21_value__36[27:17];
  assign p22_s_0__152_comb = p21_value__36[20:7] ^ p21_value__36[31:18] ^ p21_value__36[16:3];
  assign p22_temp1__398_comb = p21_e__23 + p22_S1__26_comb;
  assign p22_temp1__399_comb = p22_ch__26_comb + p22_temp1__284_comb;
  assign p22_temp2__25_comb = p22_S0__25_comb + p22_maj__25_comb;
  assign p22_value__77_comb = p21_value__57 + p22_s_1__26_comb;
  assign p22_s_0__27_comb = {p22_s_0__155_comb, p22_s_0__154_comb, p22_s_0__153_comb, p22_s_0__152_comb};
  assign p22_temp1__400_comb = p22_temp1__398_comb + p22_temp1__399_comb;
  assign p22_a__26_comb = p22_temp1__104_comb + p22_temp2__25_comb;
  assign p22_value__78_comb = p21_value__76 + p22_value__77_comb;
  assign p22_value__79_comb = p21_value__33 + p22_s_0__27_comb;

  // Registers for pipe stage 22:
  reg [31:0] p22_e__24;
  reg [31:0] p22_e__25;
  reg [31:0] p22_e__26;
  reg [31:0] p22_a__23;
  reg [31:0] p22_temp1__400;
  reg [31:0] p22_value__36;
  reg [31:0] p22_a__24;
  reg [31:0] p22_value__39;
  reg [31:0] p22_a__25;
  reg [31:0] p22_and_59596;
  reg [31:0] p22_value__42;
  reg [31:0] p22_a__26;
  reg [31:0] p22_value__45;
  reg [31:0] p22_value__48;
  reg [31:0] p22_value__51;
  reg [31:0] p22_value__54;
  reg [31:0] p22_value__57;
  reg [31:0] p22_value__60;
  reg [31:0] p22_value__61;
  reg [31:0] p22_value__66;
  reg [31:0] p22_value__67;
  reg [31:0] p22_value__72;
  reg [31:0] p22_value__73;
  reg [31:0] p22_value__78;
  reg [31:0] p22_value__79;
  always_ff @ (posedge clk) begin
    p22_e__24 <= p21_e__24;
    p22_e__25 <= p21_e__25;
    p22_e__26 <= p22_e__26_comb;
    p22_a__23 <= p21_a__23;
    p22_temp1__400 <= p22_temp1__400_comb;
    p22_value__36 <= p21_value__36;
    p22_a__24 <= p21_a__24;
    p22_value__39 <= p21_value__39;
    p22_a__25 <= p21_a__25;
    p22_and_59596 <= p22_and_59596_comb;
    p22_value__42 <= p21_value__42;
    p22_a__26 <= p22_a__26_comb;
    p22_value__45 <= p21_value__45;
    p22_value__48 <= p21_value__48;
    p22_value__51 <= p21_value__51;
    p22_value__54 <= p21_value__54;
    p22_value__57 <= p21_value__57;
    p22_value__60 <= p21_value__60;
    p22_value__61 <= p21_value__61;
    p22_value__66 <= p21_value__66;
    p22_value__67 <= p21_value__67;
    p22_value__72 <= p21_value__72;
    p22_value__73 <= p21_value__73;
    p22_value__78 <= p22_value__78_comb;
    p22_value__79 <= p22_value__79_comb;
  end

  // ===== Pipe stage 23:
  wire [31:0] p23_e__27_comb;
  wire [5:0] p23_S1__171_comb;
  wire [4:0] p23_S1__170_comb;
  wire [13:0] p23_S1__169_comb;
  wire [6:0] p23_S1__168_comb;
  wire [31:0] p23_S1__27_comb;
  wire [1:0] p23_S0__167_comb;
  wire [10:0] p23_S0__166_comb;
  wire [8:0] p23_S0__165_comb;
  wire [9:0] p23_S0__164_comb;
  wire [31:0] p23_and_59730_comb;
  wire [31:0] p23_temp1__109_comb;
  wire [31:0] p23_ch__27_comb;
  wire [31:0] p23_S0__26_comb;
  wire [31:0] p23_maj__26_comb;
  wire [2:0] p23_s_0__159_comb;
  wire [3:0] p23_s_0__158_comb;
  wire [10:0] p23_s_0__157_comb;
  wire [13:0] p23_s_0__156_comb;
  wire [31:0] p23_temp1__110_comb;
  wire [31:0] p23_temp1__285_comb;
  wire [31:0] p23_temp2__26_comb;
  wire [31:0] p23_s_0__28_comb;
  wire [31:0] p23_temp1__112_comb;
  wire [31:0] p23_a__27_comb;
  wire [31:0] p23_value__82_comb;
  assign p23_e__27_comb = p22_a__23 + p22_temp1__400;
  assign p23_S1__171_comb = p23_e__27_comb[5:0] ^ p23_e__27_comb[10:5] ^ p23_e__27_comb[24:19];
  assign p23_S1__170_comb = p23_e__27_comb[31:27] ^ p23_e__27_comb[4:0] ^ p23_e__27_comb[18:14];
  assign p23_S1__169_comb = p23_e__27_comb[26:13] ^ p23_e__27_comb[31:18] ^ p23_e__27_comb[13:0];
  assign p23_S1__168_comb = p23_e__27_comb[12:6] ^ p23_e__27_comb[17:11] ^ p23_e__27_comb[31:25];
  assign p23_S1__27_comb = {p23_S1__171_comb, p23_S1__170_comb, p23_S1__169_comb, p23_S1__168_comb};
  assign p23_S0__167_comb = p22_a__26[1:0] ^ p22_a__26[12:11] ^ p22_a__26[21:20];
  assign p23_S0__166_comb = p22_a__26[31:21] ^ p22_a__26[10:0] ^ p22_a__26[19:9];
  assign p23_S0__165_comb = p22_a__26[20:12] ^ p22_a__26[31:23] ^ p22_a__26[8:0];
  assign p23_S0__164_comb = p22_a__26[11:2] ^ p22_a__26[22:13] ^ p22_a__26[31:22];
  assign p23_and_59730_comb = p22_a__26 & p22_a__25;
  assign p23_temp1__109_comb = p22_e__24 + p23_S1__27_comb;
  assign p23_ch__27_comb = p23_e__27_comb & p22_e__26 ^ ~(p23_e__27_comb | ~p22_e__25);
  assign p23_S0__26_comb = {p23_S0__167_comb, p23_S0__166_comb, p23_S0__165_comb, p23_S0__164_comb};
  assign p23_maj__26_comb = p23_and_59730_comb ^ p22_a__26 & p22_a__24 ^ p22_and_59596;
  assign p23_s_0__159_comb = p22_value__39[6:4] ^ p22_value__39[17:15];
  assign p23_s_0__158_comb = p22_value__39[3:0] ^ p22_value__39[14:11] ^ p22_value__39[31:28];
  assign p23_s_0__157_comb = p22_value__39[31:21] ^ p22_value__39[10:0] ^ p22_value__39[27:17];
  assign p23_s_0__156_comb = p22_value__39[20:7] ^ p22_value__39[31:18] ^ p22_value__39[16:3];
  assign p23_temp1__110_comb = p23_temp1__109_comb + p23_ch__27_comb;
  assign p23_temp1__285_comb = p22_value__36 + 32'hbf59_7fc7;
  assign p23_temp2__26_comb = p23_S0__26_comb + p23_maj__26_comb;
  assign p23_s_0__28_comb = {p23_s_0__159_comb, p23_s_0__158_comb, p23_s_0__157_comb, p23_s_0__156_comb};
  assign p23_temp1__112_comb = p23_temp1__110_comb + p23_temp1__285_comb;
  assign p23_a__27_comb = p22_temp1__400 + p23_temp2__26_comb;
  assign p23_value__82_comb = p22_value__36 + p23_s_0__28_comb;

  // Registers for pipe stage 23:
  reg [31:0] p23_e__25;
  reg [31:0] p23_e__26;
  reg [31:0] p23_e__27;
  reg [31:0] p23_a__24;
  reg [31:0] p23_temp1__112;
  reg [31:0] p23_value__39;
  reg [31:0] p23_a__25;
  reg [31:0] p23_value__42;
  reg [31:0] p23_a__26;
  reg [31:0] p23_and_59730;
  reg [31:0] p23_value__45;
  reg [31:0] p23_a__27;
  reg [31:0] p23_value__48;
  reg [31:0] p23_value__51;
  reg [31:0] p23_value__54;
  reg [31:0] p23_value__57;
  reg [31:0] p23_value__60;
  reg [31:0] p23_value__61;
  reg [31:0] p23_value__66;
  reg [31:0] p23_value__67;
  reg [31:0] p23_value__72;
  reg [31:0] p23_value__73;
  reg [31:0] p23_value__78;
  reg [31:0] p23_value__79;
  reg [31:0] p23_value__82;
  always_ff @ (posedge clk) begin
    p23_e__25 <= p22_e__25;
    p23_e__26 <= p22_e__26;
    p23_e__27 <= p23_e__27_comb;
    p23_a__24 <= p22_a__24;
    p23_temp1__112 <= p23_temp1__112_comb;
    p23_value__39 <= p22_value__39;
    p23_a__25 <= p22_a__25;
    p23_value__42 <= p22_value__42;
    p23_a__26 <= p22_a__26;
    p23_and_59730 <= p23_and_59730_comb;
    p23_value__45 <= p22_value__45;
    p23_a__27 <= p23_a__27_comb;
    p23_value__48 <= p22_value__48;
    p23_value__51 <= p22_value__51;
    p23_value__54 <= p22_value__54;
    p23_value__57 <= p22_value__57;
    p23_value__60 <= p22_value__60;
    p23_value__61 <= p22_value__61;
    p23_value__66 <= p22_value__66;
    p23_value__67 <= p22_value__67;
    p23_value__72 <= p22_value__72;
    p23_value__73 <= p22_value__73;
    p23_value__78 <= p22_value__78;
    p23_value__79 <= p22_value__79;
    p23_value__82 <= p23_value__82_comb;
  end

  // ===== Pipe stage 24:
  wire [31:0] p24_e__28_comb;
  wire [5:0] p24_S1__175_comb;
  wire [4:0] p24_S1__174_comb;
  wire [13:0] p24_S1__173_comb;
  wire [6:0] p24_S1__172_comb;
  wire [31:0] p24_S1__28_comb;
  wire [1:0] p24_S0__171_comb;
  wire [10:0] p24_S0__170_comb;
  wire [8:0] p24_S0__169_comb;
  wire [9:0] p24_S0__168_comb;
  wire [31:0] p24_and_59846_comb;
  wire [31:0] p24_temp1__113_comb;
  wire [31:0] p24_ch__28_comb;
  wire [31:0] p24_S0__27_comb;
  wire [31:0] p24_maj__27_comb;
  wire [2:0] p24_s_0__163_comb;
  wire [3:0] p24_s_0__162_comb;
  wire [10:0] p24_s_0__161_comb;
  wire [13:0] p24_s_0__160_comb;
  wire [31:0] p24_temp1__114_comb;
  wire [31:0] p24_temp1__286_comb;
  wire [31:0] p24_temp2__27_comb;
  wire [31:0] p24_s_0__29_comb;
  wire [31:0] p24_temp1__116_comb;
  wire [31:0] p24_a__28_comb;
  wire [31:0] p24_value__85_comb;
  assign p24_e__28_comb = p23_a__24 + p23_temp1__112;
  assign p24_S1__175_comb = p24_e__28_comb[5:0] ^ p24_e__28_comb[10:5] ^ p24_e__28_comb[24:19];
  assign p24_S1__174_comb = p24_e__28_comb[31:27] ^ p24_e__28_comb[4:0] ^ p24_e__28_comb[18:14];
  assign p24_S1__173_comb = p24_e__28_comb[26:13] ^ p24_e__28_comb[31:18] ^ p24_e__28_comb[13:0];
  assign p24_S1__172_comb = p24_e__28_comb[12:6] ^ p24_e__28_comb[17:11] ^ p24_e__28_comb[31:25];
  assign p24_S1__28_comb = {p24_S1__175_comb, p24_S1__174_comb, p24_S1__173_comb, p24_S1__172_comb};
  assign p24_S0__171_comb = p23_a__27[1:0] ^ p23_a__27[12:11] ^ p23_a__27[21:20];
  assign p24_S0__170_comb = p23_a__27[31:21] ^ p23_a__27[10:0] ^ p23_a__27[19:9];
  assign p24_S0__169_comb = p23_a__27[20:12] ^ p23_a__27[31:23] ^ p23_a__27[8:0];
  assign p24_S0__168_comb = p23_a__27[11:2] ^ p23_a__27[22:13] ^ p23_a__27[31:22];
  assign p24_and_59846_comb = p23_a__27 & p23_a__26;
  assign p24_temp1__113_comb = p23_e__25 + p24_S1__28_comb;
  assign p24_ch__28_comb = p24_e__28_comb & p23_e__27 ^ ~(p24_e__28_comb | ~p23_e__26);
  assign p24_S0__27_comb = {p24_S0__171_comb, p24_S0__170_comb, p24_S0__169_comb, p24_S0__168_comb};
  assign p24_maj__27_comb = p24_and_59846_comb ^ p23_a__27 & p23_a__25 ^ p23_and_59730;
  assign p24_s_0__163_comb = p23_value__42[6:4] ^ p23_value__42[17:15];
  assign p24_s_0__162_comb = p23_value__42[3:0] ^ p23_value__42[14:11] ^ p23_value__42[31:28];
  assign p24_s_0__161_comb = p23_value__42[31:21] ^ p23_value__42[10:0] ^ p23_value__42[27:17];
  assign p24_s_0__160_comb = p23_value__42[20:7] ^ p23_value__42[31:18] ^ p23_value__42[16:3];
  assign p24_temp1__114_comb = p24_temp1__113_comb + p24_ch__28_comb;
  assign p24_temp1__286_comb = p23_value__39 + 32'hc6e0_0bf3;
  assign p24_temp2__27_comb = p24_S0__27_comb + p24_maj__27_comb;
  assign p24_s_0__29_comb = {p24_s_0__163_comb, p24_s_0__162_comb, p24_s_0__161_comb, p24_s_0__160_comb};
  assign p24_temp1__116_comb = p24_temp1__114_comb + p24_temp1__286_comb;
  assign p24_a__28_comb = p23_temp1__112 + p24_temp2__27_comb;
  assign p24_value__85_comb = p23_value__39 + p24_s_0__29_comb;

  // Registers for pipe stage 24:
  reg [31:0] p24_e__26;
  reg [31:0] p24_e__27;
  reg [31:0] p24_e__28;
  reg [31:0] p24_a__25;
  reg [31:0] p24_temp1__116;
  reg [31:0] p24_value__42;
  reg [31:0] p24_a__26;
  reg [31:0] p24_value__45;
  reg [31:0] p24_a__27;
  reg [31:0] p24_and_59846;
  reg [31:0] p24_value__48;
  reg [31:0] p24_a__28;
  reg [31:0] p24_value__51;
  reg [31:0] p24_value__54;
  reg [31:0] p24_value__57;
  reg [31:0] p24_value__60;
  reg [31:0] p24_value__61;
  reg [31:0] p24_value__66;
  reg [31:0] p24_value__67;
  reg [31:0] p24_value__72;
  reg [31:0] p24_value__73;
  reg [31:0] p24_value__78;
  reg [31:0] p24_value__79;
  reg [31:0] p24_value__82;
  reg [31:0] p24_value__85;
  always_ff @ (posedge clk) begin
    p24_e__26 <= p23_e__26;
    p24_e__27 <= p23_e__27;
    p24_e__28 <= p24_e__28_comb;
    p24_a__25 <= p23_a__25;
    p24_temp1__116 <= p24_temp1__116_comb;
    p24_value__42 <= p23_value__42;
    p24_a__26 <= p23_a__26;
    p24_value__45 <= p23_value__45;
    p24_a__27 <= p23_a__27;
    p24_and_59846 <= p24_and_59846_comb;
    p24_value__48 <= p23_value__48;
    p24_a__28 <= p24_a__28_comb;
    p24_value__51 <= p23_value__51;
    p24_value__54 <= p23_value__54;
    p24_value__57 <= p23_value__57;
    p24_value__60 <= p23_value__60;
    p24_value__61 <= p23_value__61;
    p24_value__66 <= p23_value__66;
    p24_value__67 <= p23_value__67;
    p24_value__72 <= p23_value__72;
    p24_value__73 <= p23_value__73;
    p24_value__78 <= p23_value__78;
    p24_value__79 <= p23_value__79;
    p24_value__82 <= p23_value__82;
    p24_value__85 <= p24_value__85_comb;
  end

  // ===== Pipe stage 25:
  wire [31:0] p25_e__29_comb;
  wire [5:0] p25_S1__179_comb;
  wire [4:0] p25_S1__178_comb;
  wire [13:0] p25_S1__177_comb;
  wire [6:0] p25_S1__176_comb;
  wire [31:0] p25_S1__29_comb;
  wire [1:0] p25_S0__175_comb;
  wire [10:0] p25_S0__174_comb;
  wire [8:0] p25_S0__173_comb;
  wire [9:0] p25_S0__172_comb;
  wire [31:0] p25_and_59962_comb;
  wire [31:0] p25_temp1__117_comb;
  wire [31:0] p25_ch__29_comb;
  wire [31:0] p25_S0__28_comb;
  wire [31:0] p25_maj__28_comb;
  wire [31:0] p25_temp1__118_comb;
  wire [31:0] p25_temp1__287_comb;
  wire [31:0] p25_temp2__28_comb;
  wire [31:0] p25_temp1__120_comb;
  wire [31:0] p25_a__29_comb;
  assign p25_e__29_comb = p24_a__25 + p24_temp1__116;
  assign p25_S1__179_comb = p25_e__29_comb[5:0] ^ p25_e__29_comb[10:5] ^ p25_e__29_comb[24:19];
  assign p25_S1__178_comb = p25_e__29_comb[31:27] ^ p25_e__29_comb[4:0] ^ p25_e__29_comb[18:14];
  assign p25_S1__177_comb = p25_e__29_comb[26:13] ^ p25_e__29_comb[31:18] ^ p25_e__29_comb[13:0];
  assign p25_S1__176_comb = p25_e__29_comb[12:6] ^ p25_e__29_comb[17:11] ^ p25_e__29_comb[31:25];
  assign p25_S1__29_comb = {p25_S1__179_comb, p25_S1__178_comb, p25_S1__177_comb, p25_S1__176_comb};
  assign p25_S0__175_comb = p24_a__28[1:0] ^ p24_a__28[12:11] ^ p24_a__28[21:20];
  assign p25_S0__174_comb = p24_a__28[31:21] ^ p24_a__28[10:0] ^ p24_a__28[19:9];
  assign p25_S0__173_comb = p24_a__28[20:12] ^ p24_a__28[31:23] ^ p24_a__28[8:0];
  assign p25_S0__172_comb = p24_a__28[11:2] ^ p24_a__28[22:13] ^ p24_a__28[31:22];
  assign p25_and_59962_comb = p24_a__28 & p24_a__27;
  assign p25_temp1__117_comb = p24_e__26 + p25_S1__29_comb;
  assign p25_ch__29_comb = p25_e__29_comb & p24_e__28 ^ ~(p25_e__29_comb | ~p24_e__27);
  assign p25_S0__28_comb = {p25_S0__175_comb, p25_S0__174_comb, p25_S0__173_comb, p25_S0__172_comb};
  assign p25_maj__28_comb = p25_and_59962_comb ^ p24_a__28 & p24_a__26 ^ p24_and_59846;
  assign p25_temp1__118_comb = p25_temp1__117_comb + p25_ch__29_comb;
  assign p25_temp1__287_comb = p24_value__42 + 32'hd5a7_9147;
  assign p25_temp2__28_comb = p25_S0__28_comb + p25_maj__28_comb;
  assign p25_temp1__120_comb = p25_temp1__118_comb + p25_temp1__287_comb;
  assign p25_a__29_comb = p24_temp1__116 + p25_temp2__28_comb;

  // Registers for pipe stage 25:
  reg [31:0] p25_e__27;
  reg [31:0] p25_e__28;
  reg [31:0] p25_e__29;
  reg [31:0] p25_value__42;
  reg [31:0] p25_a__26;
  reg [31:0] p25_temp1__120;
  reg [31:0] p25_value__45;
  reg [31:0] p25_a__27;
  reg [31:0] p25_value__48;
  reg [31:0] p25_a__28;
  reg [31:0] p25_and_59962;
  reg [31:0] p25_value__51;
  reg [31:0] p25_a__29;
  reg [31:0] p25_value__54;
  reg [31:0] p25_value__57;
  reg [31:0] p25_value__60;
  reg [31:0] p25_value__61;
  reg [31:0] p25_value__66;
  reg [31:0] p25_value__67;
  reg [31:0] p25_value__72;
  reg [31:0] p25_value__73;
  reg [31:0] p25_value__78;
  reg [31:0] p25_value__79;
  reg [31:0] p25_value__82;
  reg [31:0] p25_value__85;
  always_ff @ (posedge clk) begin
    p25_e__27 <= p24_e__27;
    p25_e__28 <= p24_e__28;
    p25_e__29 <= p25_e__29_comb;
    p25_value__42 <= p24_value__42;
    p25_a__26 <= p24_a__26;
    p25_temp1__120 <= p25_temp1__120_comb;
    p25_value__45 <= p24_value__45;
    p25_a__27 <= p24_a__27;
    p25_value__48 <= p24_value__48;
    p25_a__28 <= p24_a__28;
    p25_and_59962 <= p25_and_59962_comb;
    p25_value__51 <= p24_value__51;
    p25_a__29 <= p25_a__29_comb;
    p25_value__54 <= p24_value__54;
    p25_value__57 <= p24_value__57;
    p25_value__60 <= p24_value__60;
    p25_value__61 <= p24_value__61;
    p25_value__66 <= p24_value__66;
    p25_value__67 <= p24_value__67;
    p25_value__72 <= p24_value__72;
    p25_value__73 <= p24_value__73;
    p25_value__78 <= p24_value__78;
    p25_value__79 <= p24_value__79;
    p25_value__82 <= p24_value__82;
    p25_value__85 <= p24_value__85;
  end

  // ===== Pipe stage 26:
  wire [31:0] p26_e__30_comb;
  wire [5:0] p26_S1__183_comb;
  wire [4:0] p26_S1__182_comb;
  wire [13:0] p26_S1__181_comb;
  wire [6:0] p26_S1__180_comb;
  wire [31:0] p26_S1__30_comb;
  wire [1:0] p26_S0__179_comb;
  wire [10:0] p26_S0__178_comb;
  wire [8:0] p26_S0__177_comb;
  wire [9:0] p26_S0__176_comb;
  wire [31:0] p26_and_60061_comb;
  wire [31:0] p26_temp1__121_comb;
  wire [31:0] p26_ch__30_comb;
  wire [31:0] p26_S0__29_comb;
  wire [31:0] p26_maj__29_comb;
  wire [31:0] p26_temp1__122_comb;
  wire [31:0] p26_temp1__288_comb;
  wire [31:0] p26_temp2__29_comb;
  wire [31:0] p26_temp1__124_comb;
  wire [31:0] p26_a__30_comb;
  assign p26_e__30_comb = p25_a__26 + p25_temp1__120;
  assign p26_S1__183_comb = p26_e__30_comb[5:0] ^ p26_e__30_comb[10:5] ^ p26_e__30_comb[24:19];
  assign p26_S1__182_comb = p26_e__30_comb[31:27] ^ p26_e__30_comb[4:0] ^ p26_e__30_comb[18:14];
  assign p26_S1__181_comb = p26_e__30_comb[26:13] ^ p26_e__30_comb[31:18] ^ p26_e__30_comb[13:0];
  assign p26_S1__180_comb = p26_e__30_comb[12:6] ^ p26_e__30_comb[17:11] ^ p26_e__30_comb[31:25];
  assign p26_S1__30_comb = {p26_S1__183_comb, p26_S1__182_comb, p26_S1__181_comb, p26_S1__180_comb};
  assign p26_S0__179_comb = p25_a__29[1:0] ^ p25_a__29[12:11] ^ p25_a__29[21:20];
  assign p26_S0__178_comb = p25_a__29[31:21] ^ p25_a__29[10:0] ^ p25_a__29[19:9];
  assign p26_S0__177_comb = p25_a__29[20:12] ^ p25_a__29[31:23] ^ p25_a__29[8:0];
  assign p26_S0__176_comb = p25_a__29[11:2] ^ p25_a__29[22:13] ^ p25_a__29[31:22];
  assign p26_and_60061_comb = p25_a__29 & p25_a__28;
  assign p26_temp1__121_comb = p25_e__27 + p26_S1__30_comb;
  assign p26_ch__30_comb = p26_e__30_comb & p25_e__29 ^ ~(p26_e__30_comb | ~p25_e__28);
  assign p26_S0__29_comb = {p26_S0__179_comb, p26_S0__178_comb, p26_S0__177_comb, p26_S0__176_comb};
  assign p26_maj__29_comb = p26_and_60061_comb ^ p25_a__29 & p25_a__27 ^ p25_and_59962;
  assign p26_temp1__122_comb = p26_temp1__121_comb + p26_ch__30_comb;
  assign p26_temp1__288_comb = p25_value__45 + 32'h06ca_6351;
  assign p26_temp2__29_comb = p26_S0__29_comb + p26_maj__29_comb;
  assign p26_temp1__124_comb = p26_temp1__122_comb + p26_temp1__288_comb;
  assign p26_a__30_comb = p25_temp1__120 + p26_temp2__29_comb;

  // Registers for pipe stage 26:
  reg [31:0] p26_e__28;
  reg [31:0] p26_e__29;
  reg [31:0] p26_value__42;
  reg [31:0] p26_e__30;
  reg [31:0] p26_value__45;
  reg [31:0] p26_a__27;
  reg [31:0] p26_temp1__124;
  reg [31:0] p26_value__48;
  reg [31:0] p26_a__28;
  reg [31:0] p26_value__51;
  reg [31:0] p26_a__29;
  reg [31:0] p26_value__54;
  reg [31:0] p26_and_60061;
  reg [31:0] p26_a__30;
  reg [31:0] p26_value__57;
  reg [31:0] p26_value__60;
  reg [31:0] p26_value__61;
  reg [31:0] p26_value__66;
  reg [31:0] p26_value__67;
  reg [31:0] p26_value__72;
  reg [31:0] p26_value__73;
  reg [31:0] p26_value__78;
  reg [31:0] p26_value__79;
  reg [31:0] p26_value__82;
  reg [31:0] p26_value__85;
  always_ff @ (posedge clk) begin
    p26_e__28 <= p25_e__28;
    p26_e__29 <= p25_e__29;
    p26_value__42 <= p25_value__42;
    p26_e__30 <= p26_e__30_comb;
    p26_value__45 <= p25_value__45;
    p26_a__27 <= p25_a__27;
    p26_temp1__124 <= p26_temp1__124_comb;
    p26_value__48 <= p25_value__48;
    p26_a__28 <= p25_a__28;
    p26_value__51 <= p25_value__51;
    p26_a__29 <= p25_a__29;
    p26_value__54 <= p25_value__54;
    p26_and_60061 <= p26_and_60061_comb;
    p26_a__30 <= p26_a__30_comb;
    p26_value__57 <= p25_value__57;
    p26_value__60 <= p25_value__60;
    p26_value__61 <= p25_value__61;
    p26_value__66 <= p25_value__66;
    p26_value__67 <= p25_value__67;
    p26_value__72 <= p25_value__72;
    p26_value__73 <= p25_value__73;
    p26_value__78 <= p25_value__78;
    p26_value__79 <= p25_value__79;
    p26_value__82 <= p25_value__82;
    p26_value__85 <= p25_value__85;
  end

  // ===== Pipe stage 27:
  wire [31:0] p27_e__31_comb;
  wire [5:0] p27_S1__187_comb;
  wire [4:0] p27_S1__186_comb;
  wire [13:0] p27_S1__185_comb;
  wire [6:0] p27_S1__184_comb;
  wire [31:0] p27_S1__31_comb;
  wire [1:0] p27_S0__183_comb;
  wire [10:0] p27_S0__182_comb;
  wire [8:0] p27_S0__181_comb;
  wire [9:0] p27_S0__180_comb;
  wire [31:0] p27_and_60160_comb;
  wire [31:0] p27_temp1__125_comb;
  wire [31:0] p27_ch__31_comb;
  wire [31:0] p27_S0__30_comb;
  wire [31:0] p27_maj__30_comb;
  wire [31:0] p27_temp1__126_comb;
  wire [31:0] p27_temp1__289_comb;
  wire [31:0] p27_temp2__30_comb;
  wire [31:0] p27_temp1__128_comb;
  wire [31:0] p27_a__31_comb;
  assign p27_e__31_comb = p26_a__27 + p26_temp1__124;
  assign p27_S1__187_comb = p27_e__31_comb[5:0] ^ p27_e__31_comb[10:5] ^ p27_e__31_comb[24:19];
  assign p27_S1__186_comb = p27_e__31_comb[31:27] ^ p27_e__31_comb[4:0] ^ p27_e__31_comb[18:14];
  assign p27_S1__185_comb = p27_e__31_comb[26:13] ^ p27_e__31_comb[31:18] ^ p27_e__31_comb[13:0];
  assign p27_S1__184_comb = p27_e__31_comb[12:6] ^ p27_e__31_comb[17:11] ^ p27_e__31_comb[31:25];
  assign p27_S1__31_comb = {p27_S1__187_comb, p27_S1__186_comb, p27_S1__185_comb, p27_S1__184_comb};
  assign p27_S0__183_comb = p26_a__30[1:0] ^ p26_a__30[12:11] ^ p26_a__30[21:20];
  assign p27_S0__182_comb = p26_a__30[31:21] ^ p26_a__30[10:0] ^ p26_a__30[19:9];
  assign p27_S0__181_comb = p26_a__30[20:12] ^ p26_a__30[31:23] ^ p26_a__30[8:0];
  assign p27_S0__180_comb = p26_a__30[11:2] ^ p26_a__30[22:13] ^ p26_a__30[31:22];
  assign p27_and_60160_comb = p26_a__30 & p26_a__29;
  assign p27_temp1__125_comb = p26_e__28 + p27_S1__31_comb;
  assign p27_ch__31_comb = p27_e__31_comb & p26_e__30 ^ ~(p27_e__31_comb | ~p26_e__29);
  assign p27_S0__30_comb = {p27_S0__183_comb, p27_S0__182_comb, p27_S0__181_comb, p27_S0__180_comb};
  assign p27_maj__30_comb = p27_and_60160_comb ^ p26_a__30 & p26_a__28 ^ p26_and_60061;
  assign p27_temp1__126_comb = p27_temp1__125_comb + p27_ch__31_comb;
  assign p27_temp1__289_comb = p26_value__48 + 32'h1429_2967;
  assign p27_temp2__30_comb = p27_S0__30_comb + p27_maj__30_comb;
  assign p27_temp1__128_comb = p27_temp1__126_comb + p27_temp1__289_comb;
  assign p27_a__31_comb = p26_temp1__124 + p27_temp2__30_comb;

  // Registers for pipe stage 27:
  reg [31:0] p27_e__29;
  reg [31:0] p27_value__42;
  reg [31:0] p27_e__30;
  reg [31:0] p27_value__45;
  reg [31:0] p27_e__31;
  reg [31:0] p27_value__48;
  reg [31:0] p27_a__28;
  reg [31:0] p27_temp1__128;
  reg [31:0] p27_value__51;
  reg [31:0] p27_a__29;
  reg [31:0] p27_value__54;
  reg [31:0] p27_a__30;
  reg [31:0] p27_value__57;
  reg [31:0] p27_and_60160;
  reg [31:0] p27_a__31;
  reg [31:0] p27_value__60;
  reg [31:0] p27_value__61;
  reg [31:0] p27_value__66;
  reg [31:0] p27_value__67;
  reg [31:0] p27_value__72;
  reg [31:0] p27_value__73;
  reg [31:0] p27_value__78;
  reg [31:0] p27_value__79;
  reg [31:0] p27_value__82;
  reg [31:0] p27_value__85;
  always_ff @ (posedge clk) begin
    p27_e__29 <= p26_e__29;
    p27_value__42 <= p26_value__42;
    p27_e__30 <= p26_e__30;
    p27_value__45 <= p26_value__45;
    p27_e__31 <= p27_e__31_comb;
    p27_value__48 <= p26_value__48;
    p27_a__28 <= p26_a__28;
    p27_temp1__128 <= p27_temp1__128_comb;
    p27_value__51 <= p26_value__51;
    p27_a__29 <= p26_a__29;
    p27_value__54 <= p26_value__54;
    p27_a__30 <= p26_a__30;
    p27_value__57 <= p26_value__57;
    p27_and_60160 <= p27_and_60160_comb;
    p27_a__31 <= p27_a__31_comb;
    p27_value__60 <= p26_value__60;
    p27_value__61 <= p26_value__61;
    p27_value__66 <= p26_value__66;
    p27_value__67 <= p26_value__67;
    p27_value__72 <= p26_value__72;
    p27_value__73 <= p26_value__73;
    p27_value__78 <= p26_value__78;
    p27_value__79 <= p26_value__79;
    p27_value__82 <= p26_value__82;
    p27_value__85 <= p26_value__85;
  end

  // ===== Pipe stage 28:
  wire [31:0] p28_e__32_comb;
  wire [5:0] p28_S1__191_comb;
  wire [4:0] p28_S1__190_comb;
  wire [13:0] p28_S1__189_comb;
  wire [6:0] p28_S1__188_comb;
  wire [31:0] p28_S1__32_comb;
  wire [1:0] p28_S0__187_comb;
  wire [10:0] p28_S0__186_comb;
  wire [8:0] p28_S0__185_comb;
  wire [9:0] p28_S0__184_comb;
  wire [31:0] p28_and_60259_comb;
  wire [31:0] p28_temp1__129_comb;
  wire [31:0] p28_ch__32_comb;
  wire [31:0] p28_S0__31_comb;
  wire [31:0] p28_maj__31_comb;
  wire [31:0] p28_temp1__130_comb;
  wire [31:0] p28_temp1__290_comb;
  wire [31:0] p28_temp2__31_comb;
  wire [31:0] p28_temp1__132_comb;
  wire [31:0] p28_a__32_comb;
  assign p28_e__32_comb = p27_a__28 + p27_temp1__128;
  assign p28_S1__191_comb = p28_e__32_comb[5:0] ^ p28_e__32_comb[10:5] ^ p28_e__32_comb[24:19];
  assign p28_S1__190_comb = p28_e__32_comb[31:27] ^ p28_e__32_comb[4:0] ^ p28_e__32_comb[18:14];
  assign p28_S1__189_comb = p28_e__32_comb[26:13] ^ p28_e__32_comb[31:18] ^ p28_e__32_comb[13:0];
  assign p28_S1__188_comb = p28_e__32_comb[12:6] ^ p28_e__32_comb[17:11] ^ p28_e__32_comb[31:25];
  assign p28_S1__32_comb = {p28_S1__191_comb, p28_S1__190_comb, p28_S1__189_comb, p28_S1__188_comb};
  assign p28_S0__187_comb = p27_a__31[1:0] ^ p27_a__31[12:11] ^ p27_a__31[21:20];
  assign p28_S0__186_comb = p27_a__31[31:21] ^ p27_a__31[10:0] ^ p27_a__31[19:9];
  assign p28_S0__185_comb = p27_a__31[20:12] ^ p27_a__31[31:23] ^ p27_a__31[8:0];
  assign p28_S0__184_comb = p27_a__31[11:2] ^ p27_a__31[22:13] ^ p27_a__31[31:22];
  assign p28_and_60259_comb = p27_a__31 & p27_a__30;
  assign p28_temp1__129_comb = p27_e__29 + p28_S1__32_comb;
  assign p28_ch__32_comb = p28_e__32_comb & p27_e__31 ^ ~(p28_e__32_comb | ~p27_e__30);
  assign p28_S0__31_comb = {p28_S0__187_comb, p28_S0__186_comb, p28_S0__185_comb, p28_S0__184_comb};
  assign p28_maj__31_comb = p28_and_60259_comb ^ p27_a__31 & p27_a__29 ^ p27_and_60160;
  assign p28_temp1__130_comb = p28_temp1__129_comb + p28_ch__32_comb;
  assign p28_temp1__290_comb = p27_value__51 + 32'h27b7_0a85;
  assign p28_temp2__31_comb = p28_S0__31_comb + p28_maj__31_comb;
  assign p28_temp1__132_comb = p28_temp1__130_comb + p28_temp1__290_comb;
  assign p28_a__32_comb = p27_temp1__128 + p28_temp2__31_comb;

  // Registers for pipe stage 28:
  reg [31:0] p28_value__42;
  reg [31:0] p28_e__30;
  reg [31:0] p28_value__45;
  reg [31:0] p28_e__31;
  reg [31:0] p28_value__48;
  reg [31:0] p28_e__32;
  reg [31:0] p28_value__51;
  reg [31:0] p28_a__29;
  reg [31:0] p28_temp1__132;
  reg [31:0] p28_value__54;
  reg [31:0] p28_a__30;
  reg [31:0] p28_value__57;
  reg [31:0] p28_a__31;
  reg [31:0] p28_and_60259;
  reg [31:0] p28_value__60;
  reg [31:0] p28_a__32;
  reg [31:0] p28_value__61;
  reg [31:0] p28_value__66;
  reg [31:0] p28_value__67;
  reg [31:0] p28_value__72;
  reg [31:0] p28_value__73;
  reg [31:0] p28_value__78;
  reg [31:0] p28_value__79;
  reg [31:0] p28_value__82;
  reg [31:0] p28_value__85;
  always_ff @ (posedge clk) begin
    p28_value__42 <= p27_value__42;
    p28_e__30 <= p27_e__30;
    p28_value__45 <= p27_value__45;
    p28_e__31 <= p27_e__31;
    p28_value__48 <= p27_value__48;
    p28_e__32 <= p28_e__32_comb;
    p28_value__51 <= p27_value__51;
    p28_a__29 <= p27_a__29;
    p28_temp1__132 <= p28_temp1__132_comb;
    p28_value__54 <= p27_value__54;
    p28_a__30 <= p27_a__30;
    p28_value__57 <= p27_value__57;
    p28_a__31 <= p27_a__31;
    p28_and_60259 <= p28_and_60259_comb;
    p28_value__60 <= p27_value__60;
    p28_a__32 <= p28_a__32_comb;
    p28_value__61 <= p27_value__61;
    p28_value__66 <= p27_value__66;
    p28_value__67 <= p27_value__67;
    p28_value__72 <= p27_value__72;
    p28_value__73 <= p27_value__73;
    p28_value__78 <= p27_value__78;
    p28_value__79 <= p27_value__79;
    p28_value__82 <= p27_value__82;
    p28_value__85 <= p27_value__85;
  end

  // ===== Pipe stage 29:
  wire [1:0] p29_S0__191_comb;
  wire [10:0] p29_S0__190_comb;
  wire [8:0] p29_S0__189_comb;
  wire [9:0] p29_S0__188_comb;
  wire [31:0] p29_and_60365_comb;
  wire [31:0] p29_S0__32_comb;
  wire [31:0] p29_maj__32_comb;
  wire [31:0] p29_e__33_comb;
  wire [31:0] p29_temp2__32_comb;
  wire [31:0] p29_a__33_comb;
  wire [5:0] p29_S1__195_comb;
  wire [4:0] p29_S1__194_comb;
  wire [13:0] p29_S1__193_comb;
  wire [6:0] p29_S1__192_comb;
  wire [28:0] p29_add_60337_comb;
  wire [31:0] p29_S1__33_comb;
  wire [31:0] p29_ch__33_comb;
  wire [31:0] p29_temp1__291_comb;
  wire [1:0] p29_S0__195_comb;
  wire [10:0] p29_S0__194_comb;
  wire [8:0] p29_S0__193_comb;
  wire [9:0] p29_S0__192_comb;
  wire [31:0] p29_and_60387_comb;
  wire [31:0] p29_temp1__395_comb;
  wire [31:0] p29_temp1__396_comb;
  wire [31:0] p29_S0__33_comb;
  wire [31:0] p29_maj__33_comb;
  wire [31:0] p29_temp1__397_comb;
  wire [31:0] p29_temp2__33_comb;
  wire [31:0] p29_e__34_comb;
  wire [29:0] p29_add_60348_comb;
  wire [31:0] p29_a__34_comb;
  assign p29_S0__191_comb = p28_a__32[1:0] ^ p28_a__32[12:11] ^ p28_a__32[21:20];
  assign p29_S0__190_comb = p28_a__32[31:21] ^ p28_a__32[10:0] ^ p28_a__32[19:9];
  assign p29_S0__189_comb = p28_a__32[20:12] ^ p28_a__32[31:23] ^ p28_a__32[8:0];
  assign p29_S0__188_comb = p28_a__32[11:2] ^ p28_a__32[22:13] ^ p28_a__32[31:22];
  assign p29_and_60365_comb = p28_a__32 & p28_a__31;
  assign p29_S0__32_comb = {p29_S0__191_comb, p29_S0__190_comb, p29_S0__189_comb, p29_S0__188_comb};
  assign p29_maj__32_comb = p29_and_60365_comb ^ p28_a__32 & p28_a__30 ^ p28_and_60259;
  assign p29_e__33_comb = p28_a__29 + p28_temp1__132;
  assign p29_temp2__32_comb = p29_S0__32_comb + p29_maj__32_comb;
  assign p29_a__33_comb = p28_temp1__132 + p29_temp2__32_comb;
  assign p29_S1__195_comb = p29_e__33_comb[5:0] ^ p29_e__33_comb[10:5] ^ p29_e__33_comb[24:19];
  assign p29_S1__194_comb = p29_e__33_comb[31:27] ^ p29_e__33_comb[4:0] ^ p29_e__33_comb[18:14];
  assign p29_S1__193_comb = p29_e__33_comb[26:13] ^ p29_e__33_comb[31:18] ^ p29_e__33_comb[13:0];
  assign p29_S1__192_comb = p29_e__33_comb[12:6] ^ p29_e__33_comb[17:11] ^ p29_e__33_comb[31:25];
  assign p29_add_60337_comb = p28_value__54[31:3] + 29'h05c3_6427;
  assign p29_S1__33_comb = {p29_S1__195_comb, p29_S1__194_comb, p29_S1__193_comb, p29_S1__192_comb};
  assign p29_ch__33_comb = p29_e__33_comb & p28_e__32 ^ ~(p29_e__33_comb | ~p28_e__31);
  assign p29_temp1__291_comb = {p29_add_60337_comb, p28_value__54[2:0]};
  assign p29_S0__195_comb = p29_a__33_comb[1:0] ^ p29_a__33_comb[12:11] ^ p29_a__33_comb[21:20];
  assign p29_S0__194_comb = p29_a__33_comb[31:21] ^ p29_a__33_comb[10:0] ^ p29_a__33_comb[19:9];
  assign p29_S0__193_comb = p29_a__33_comb[20:12] ^ p29_a__33_comb[31:23] ^ p29_a__33_comb[8:0];
  assign p29_S0__192_comb = p29_a__33_comb[11:2] ^ p29_a__33_comb[22:13] ^ p29_a__33_comb[31:22];
  assign p29_and_60387_comb = p29_a__33_comb & p28_a__32;
  assign p29_temp1__395_comb = p28_e__30 + p29_S1__33_comb;
  assign p29_temp1__396_comb = p29_ch__33_comb + p29_temp1__291_comb;
  assign p29_S0__33_comb = {p29_S0__195_comb, p29_S0__194_comb, p29_S0__193_comb, p29_S0__192_comb};
  assign p29_maj__33_comb = p29_and_60387_comb ^ p29_a__33_comb & p28_a__31 ^ p29_and_60365_comb;
  assign p29_temp1__397_comb = p29_temp1__395_comb + p29_temp1__396_comb;
  assign p29_temp2__33_comb = p29_S0__33_comb + p29_maj__33_comb;
  assign p29_e__34_comb = p28_a__30 + p29_temp1__397_comb;
  assign p29_add_60348_comb = p28_value__57[31:2] + 30'h134b_1b7f;
  assign p29_a__34_comb = p29_temp1__397_comb + p29_temp2__33_comb;

  // Registers for pipe stage 29:
  reg [31:0] p29_value__42;
  reg [31:0] p29_value__45;
  reg [31:0] p29_e__31;
  reg [31:0] p29_value__48;
  reg [31:0] p29_e__32;
  reg [31:0] p29_value__51;
  reg [31:0] p29_e__33;
  reg [31:0] p29_value__54;
  reg [31:0] p29_e__34;
  reg [31:0] p29_value__57;
  reg [29:0] p29_add_60348;
  reg [31:0] p29_a__31;
  reg [31:0] p29_value__60;
  reg [31:0] p29_a__32;
  reg [31:0] p29_value__61;
  reg [31:0] p29_a__33;
  reg [31:0] p29_and_60387;
  reg [31:0] p29_value__66;
  reg [31:0] p29_a__34;
  reg [31:0] p29_value__67;
  reg [31:0] p29_value__72;
  reg [31:0] p29_value__73;
  reg [31:0] p29_value__78;
  reg [31:0] p29_value__79;
  reg [31:0] p29_value__82;
  reg [31:0] p29_value__85;
  always_ff @ (posedge clk) begin
    p29_value__42 <= p28_value__42;
    p29_value__45 <= p28_value__45;
    p29_e__31 <= p28_e__31;
    p29_value__48 <= p28_value__48;
    p29_e__32 <= p28_e__32;
    p29_value__51 <= p28_value__51;
    p29_e__33 <= p29_e__33_comb;
    p29_value__54 <= p28_value__54;
    p29_e__34 <= p29_e__34_comb;
    p29_value__57 <= p28_value__57;
    p29_add_60348 <= p29_add_60348_comb;
    p29_a__31 <= p28_a__31;
    p29_value__60 <= p28_value__60;
    p29_a__32 <= p28_a__32;
    p29_value__61 <= p28_value__61;
    p29_a__33 <= p29_a__33_comb;
    p29_and_60387 <= p29_and_60387_comb;
    p29_value__66 <= p28_value__66;
    p29_a__34 <= p29_a__34_comb;
    p29_value__67 <= p28_value__67;
    p29_value__72 <= p28_value__72;
    p29_value__73 <= p28_value__73;
    p29_value__78 <= p28_value__78;
    p29_value__79 <= p28_value__79;
    p29_value__82 <= p28_value__82;
    p29_value__85 <= p28_value__85;
  end

  // ===== Pipe stage 30:
  wire [5:0] p30_S1__199_comb;
  wire [4:0] p30_S1__198_comb;
  wire [13:0] p30_S1__197_comb;
  wire [6:0] p30_S1__196_comb;
  wire [31:0] p30_S1__34_comb;
  wire [31:0] p30_ch__34_comb;
  wire [31:0] p30_temp1__292_comb;
  wire [31:0] p30_temp1__392_comb;
  wire [31:0] p30_temp1__393_comb;
  wire [31:0] p30_temp1__394_comb;
  wire [9:0] p30_s_1__131_comb;
  wire [6:0] p30_s_1__130_comb;
  wire [1:0] p30_s_1__129_comb;
  wire [12:0] p30_s_1__128_comb;
  wire [31:0] p30_e__35_comb;
  wire [31:0] p30_s_1__21_comb;
  wire [1:0] p30_S0__199_comb;
  wire [10:0] p30_S0__198_comb;
  wire [8:0] p30_S0__197_comb;
  wire [9:0] p30_S0__196_comb;
  wire [31:0] p30_and_60523_comb;
  wire [31:0] p30_value__62_comb;
  wire [9:0] p30_s_1__159_comb;
  wire [6:0] p30_s_1__158_comb;
  wire [1:0] p30_s_1__157_comb;
  wire [12:0] p30_s_1__156_comb;
  wire [5:0] p30_S1__203_comb;
  wire [4:0] p30_S1__202_comb;
  wire [13:0] p30_S1__201_comb;
  wire [6:0] p30_S1__200_comb;
  wire [31:0] p30_S0__34_comb;
  wire [31:0] p30_maj__34_comb;
  wire [31:0] p30_value__63_comb;
  wire [31:0] p30_s_1__28_comb;
  wire [2:0] p30_s_0__167_comb;
  wire [3:0] p30_s_0__166_comb;
  wire [10:0] p30_s_0__165_comb;
  wire [13:0] p30_s_0__164_comb;
  wire [2:0] p30_s_0__171_comb;
  wire [3:0] p30_s_0__170_comb;
  wire [10:0] p30_s_0__169_comb;
  wire [13:0] p30_s_0__168_comb;
  wire [31:0] p30_S1__35_comb;
  wire [31:0] p30_temp2__34_comb;
  wire [31:0] p30_value__83_comb;
  wire [31:0] p30_s_0__30_comb;
  wire [31:0] p30_s_0__31_comb;
  wire [31:0] p30_temp1__141_comb;
  wire [31:0] p30_a__35_comb;
  wire [31:0] p30_value__84_comb;
  wire [31:0] p30_value__88_comb;
  wire [31:0] p30_value__91_comb;
  assign p30_S1__199_comb = p29_e__34[5:0] ^ p29_e__34[10:5] ^ p29_e__34[24:19];
  assign p30_S1__198_comb = p29_e__34[31:27] ^ p29_e__34[4:0] ^ p29_e__34[18:14];
  assign p30_S1__197_comb = p29_e__34[26:13] ^ p29_e__34[31:18] ^ p29_e__34[13:0];
  assign p30_S1__196_comb = p29_e__34[12:6] ^ p29_e__34[17:11] ^ p29_e__34[31:25];
  assign p30_S1__34_comb = {p30_S1__199_comb, p30_S1__198_comb, p30_S1__197_comb, p30_S1__196_comb};
  assign p30_ch__34_comb = p29_e__34 & p29_e__33 ^ ~(p29_e__34 | ~p29_e__32);
  assign p30_temp1__292_comb = {p29_add_60348, p29_value__57[1:0]};
  assign p30_temp1__392_comb = p29_e__31 + p30_S1__34_comb;
  assign p30_temp1__393_comb = p30_ch__34_comb + p30_temp1__292_comb;
  assign p30_temp1__394_comb = p30_temp1__392_comb + p30_temp1__393_comb;
  assign p30_s_1__131_comb = p29_value__57[16:7] ^ p29_value__57[18:9];
  assign p30_s_1__130_comb = p29_value__57[6:0] ^ p29_value__57[8:2] ^ p29_value__57[31:25];
  assign p30_s_1__129_comb = p29_value__57[31:30] ^ p29_value__57[1:0] ^ p29_value__57[24:23];
  assign p30_s_1__128_comb = p29_value__57[29:17] ^ p29_value__57[31:19] ^ p29_value__57[22:10];
  assign p30_e__35_comb = p29_a__31 + p30_temp1__394_comb;
  assign p30_s_1__21_comb = {p30_s_1__131_comb, p30_s_1__130_comb, p30_s_1__129_comb, p30_s_1__128_comb};
  assign p30_S0__199_comb = p29_a__34[1:0] ^ p29_a__34[12:11] ^ p29_a__34[21:20];
  assign p30_S0__198_comb = p29_a__34[31:21] ^ p29_a__34[10:0] ^ p29_a__34[19:9];
  assign p30_S0__197_comb = p29_a__34[20:12] ^ p29_a__34[31:23] ^ p29_a__34[8:0];
  assign p30_S0__196_comb = p29_a__34[11:2] ^ p29_a__34[22:13] ^ p29_a__34[31:22];
  assign p30_and_60523_comb = p29_a__34 & p29_a__33;
  assign p30_value__62_comb = p29_value__42 + p30_s_1__21_comb;
  assign p30_s_1__159_comb = p29_value__78[16:7] ^ p29_value__78[18:9];
  assign p30_s_1__158_comb = p29_value__78[6:0] ^ p29_value__78[8:2] ^ p29_value__78[31:25];
  assign p30_s_1__157_comb = p29_value__78[31:30] ^ p29_value__78[1:0] ^ p29_value__78[24:23];
  assign p30_s_1__156_comb = p29_value__78[29:17] ^ p29_value__78[31:19] ^ p29_value__78[22:10];
  assign p30_S1__203_comb = p30_e__35_comb[5:0] ^ p30_e__35_comb[10:5] ^ p30_e__35_comb[24:19];
  assign p30_S1__202_comb = p30_e__35_comb[31:27] ^ p30_e__35_comb[4:0] ^ p30_e__35_comb[18:14];
  assign p30_S1__201_comb = p30_e__35_comb[26:13] ^ p30_e__35_comb[31:18] ^ p30_e__35_comb[13:0];
  assign p30_S1__200_comb = p30_e__35_comb[12:6] ^ p30_e__35_comb[17:11] ^ p30_e__35_comb[31:25];
  assign p30_S0__34_comb = {p30_S0__199_comb, p30_S0__198_comb, p30_S0__197_comb, p30_S0__196_comb};
  assign p30_maj__34_comb = p30_and_60523_comb ^ p29_a__34 & p29_a__32 ^ p29_and_60387;
  assign p30_value__63_comb = p29_value__61 + p30_value__62_comb;
  assign p30_s_1__28_comb = {p30_s_1__159_comb, p30_s_1__158_comb, p30_s_1__157_comb, p30_s_1__156_comb};
  assign p30_s_0__167_comb = p29_value__45[6:4] ^ p29_value__45[17:15];
  assign p30_s_0__166_comb = p29_value__45[3:0] ^ p29_value__45[14:11] ^ p29_value__45[31:28];
  assign p30_s_0__165_comb = p29_value__45[31:21] ^ p29_value__45[10:0] ^ p29_value__45[27:17];
  assign p30_s_0__164_comb = p29_value__45[20:7] ^ p29_value__45[31:18] ^ p29_value__45[16:3];
  assign p30_s_0__171_comb = p29_value__48[6:4] ^ p29_value__48[17:15];
  assign p30_s_0__170_comb = p29_value__48[3:0] ^ p29_value__48[14:11] ^ p29_value__48[31:28];
  assign p30_s_0__169_comb = p29_value__48[31:21] ^ p29_value__48[10:0] ^ p29_value__48[27:17];
  assign p30_s_0__168_comb = p29_value__48[20:7] ^ p29_value__48[31:18] ^ p29_value__48[16:3];
  assign p30_S1__35_comb = {p30_S1__203_comb, p30_S1__202_comb, p30_S1__201_comb, p30_S1__200_comb};
  assign p30_temp2__34_comb = p30_S0__34_comb + p30_maj__34_comb;
  assign p30_value__83_comb = p30_value__63_comb + p30_s_1__28_comb;
  assign p30_s_0__30_comb = {p30_s_0__167_comb, p30_s_0__166_comb, p30_s_0__165_comb, p30_s_0__164_comb};
  assign p30_s_0__31_comb = {p30_s_0__171_comb, p30_s_0__170_comb, p30_s_0__169_comb, p30_s_0__168_comb};
  assign p30_temp1__141_comb = p29_e__32 + p30_S1__35_comb;
  assign p30_a__35_comb = p30_temp1__394_comb + p30_temp2__34_comb;
  assign p30_value__84_comb = p29_value__82 + p30_value__83_comb;
  assign p30_value__88_comb = p29_value__42 + p30_s_0__30_comb;
  assign p30_value__91_comb = p29_value__45 + p30_s_0__31_comb;

  // Registers for pipe stage 30:
  reg [31:0] p30_value__48;
  reg [31:0] p30_value__51;
  reg [31:0] p30_e__33;
  reg [31:0] p30_value__54;
  reg [31:0] p30_e__34;
  reg [31:0] p30_value__57;
  reg [31:0] p30_e__35;
  reg [31:0] p30_temp1__141;
  reg [31:0] p30_value__60;
  reg [31:0] p30_a__32;
  reg [31:0] p30_value__63;
  reg [31:0] p30_a__33;
  reg [31:0] p30_value__66;
  reg [31:0] p30_a__34;
  reg [31:0] p30_value__67;
  reg [31:0] p30_and_60523;
  reg [31:0] p30_a__35;
  reg [31:0] p30_value__72;
  reg [31:0] p30_value__73;
  reg [31:0] p30_value__78;
  reg [31:0] p30_value__79;
  reg [31:0] p30_value__84;
  reg [31:0] p30_value__85;
  reg [31:0] p30_value__88;
  reg [31:0] p30_value__91;
  always_ff @ (posedge clk) begin
    p30_value__48 <= p29_value__48;
    p30_value__51 <= p29_value__51;
    p30_e__33 <= p29_e__33;
    p30_value__54 <= p29_value__54;
    p30_e__34 <= p29_e__34;
    p30_value__57 <= p29_value__57;
    p30_e__35 <= p30_e__35_comb;
    p30_temp1__141 <= p30_temp1__141_comb;
    p30_value__60 <= p29_value__60;
    p30_a__32 <= p29_a__32;
    p30_value__63 <= p30_value__63_comb;
    p30_a__33 <= p29_a__33;
    p30_value__66 <= p29_value__66;
    p30_a__34 <= p29_a__34;
    p30_value__67 <= p29_value__67;
    p30_and_60523 <= p30_and_60523_comb;
    p30_a__35 <= p30_a__35_comb;
    p30_value__72 <= p29_value__72;
    p30_value__73 <= p29_value__73;
    p30_value__78 <= p29_value__78;
    p30_value__79 <= p29_value__79;
    p30_value__84 <= p30_value__84_comb;
    p30_value__85 <= p29_value__85;
    p30_value__88 <= p30_value__88_comb;
    p30_value__91 <= p30_value__91_comb;
  end

  // ===== Pipe stage 31:
  wire [9:0] p31_s_1__139_comb;
  wire [6:0] p31_s_1__138_comb;
  wire [1:0] p31_s_1__137_comb;
  wire [12:0] p31_s_1__136_comb;
  wire [31:0] p31_ch__35_comb;
  wire [31:0] p31_s_1__23_comb;
  wire [31:0] p31_temp1__142_comb;
  wire [31:0] p31_temp1__293_comb;
  wire [31:0] p31_value__68_comb;
  wire [31:0] p31_temp1__144_comb;
  wire [31:0] p31_value__69_comb;
  wire [31:0] p31_e__36_comb;
  wire [1:0] p31_S0__203_comb;
  wire [10:0] p31_S0__202_comb;
  wire [8:0] p31_S0__201_comb;
  wire [9:0] p31_S0__200_comb;
  wire [31:0] p31_and_60701_comb;
  wire [9:0] p31_s_1__147_comb;
  wire [6:0] p31_s_1__146_comb;
  wire [1:0] p31_s_1__145_comb;
  wire [12:0] p31_s_1__144_comb;
  wire [9:0] p31_s_1__167_comb;
  wire [6:0] p31_s_1__166_comb;
  wire [1:0] p31_s_1__165_comb;
  wire [12:0] p31_s_1__164_comb;
  wire [5:0] p31_S1__207_comb;
  wire [4:0] p31_S1__206_comb;
  wire [13:0] p31_S1__205_comb;
  wire [6:0] p31_S1__204_comb;
  wire [29:0] p31_add_60661_comb;
  wire [31:0] p31_S0__35_comb;
  wire [31:0] p31_maj__35_comb;
  wire [31:0] p31_s_1__25_comb;
  wire [31:0] p31_s_1__30_comb;
  wire [2:0] p31_s_0__175_comb;
  wire [3:0] p31_s_0__174_comb;
  wire [10:0] p31_s_0__173_comb;
  wire [13:0] p31_s_0__172_comb;
  wire [2:0] p31_s_0__179_comb;
  wire [3:0] p31_s_0__178_comb;
  wire [10:0] p31_s_0__177_comb;
  wire [13:0] p31_s_0__176_comb;
  wire [2:0] p31_s_0__183_comb;
  wire [3:0] p31_s_0__182_comb;
  wire [10:0] p31_s_0__181_comb;
  wire [13:0] p31_s_0__180_comb;
  wire [2:0] p31_s_0__187_comb;
  wire [3:0] p31_s_0__186_comb;
  wire [10:0] p31_s_0__185_comb;
  wire [13:0] p31_s_0__184_comb;
  wire [31:0] p31_S1__36_comb;
  wire [31:0] p31_ch__36_comb;
  wire [31:0] p31_temp1__294_comb;
  wire [31:0] p31_temp2__35_comb;
  wire [31:0] p31_value__74_comb;
  wire [31:0] p31_value__89_comb;
  wire [31:0] p31_s_0__32_comb;
  wire [31:0] p31_s_0__33_comb;
  wire [31:0] p31_s_0__34_comb;
  wire [31:0] p31_s_0__35_comb;
  wire [31:0] p31_temp1__389_comb;
  wire [31:0] p31_temp1__390_comb;
  wire [31:0] p31_a__36_comb;
  wire [31:0] p31_value__75_comb;
  wire [31:0] p31_value__90_comb;
  wire [31:0] p31_value__94_comb;
  wire [31:0] p31_value__97_comb;
  wire [31:0] p31_value__100_comb;
  wire [31:0] p31_value__103_comb;
  assign p31_s_1__139_comb = p30_value__63[16:7] ^ p30_value__63[18:9];
  assign p31_s_1__138_comb = p30_value__63[6:0] ^ p30_value__63[8:2] ^ p30_value__63[31:25];
  assign p31_s_1__137_comb = p30_value__63[31:30] ^ p30_value__63[1:0] ^ p30_value__63[24:23];
  assign p31_s_1__136_comb = p30_value__63[29:17] ^ p30_value__63[31:19] ^ p30_value__63[22:10];
  assign p31_ch__35_comb = p30_e__35 & p30_e__34 ^ ~(p30_e__35 | ~p30_e__33);
  assign p31_s_1__23_comb = {p31_s_1__139_comb, p31_s_1__138_comb, p31_s_1__137_comb, p31_s_1__136_comb};
  assign p31_temp1__142_comb = p30_temp1__141 + p31_ch__35_comb;
  assign p31_temp1__293_comb = p30_value__60 + 32'h5338_0d13;
  assign p31_value__68_comb = p30_value__48 + p31_s_1__23_comb;
  assign p31_temp1__144_comb = p31_temp1__142_comb + p31_temp1__293_comb;
  assign p31_value__69_comb = p30_value__67 + p31_value__68_comb;
  assign p31_e__36_comb = p30_a__32 + p31_temp1__144_comb;
  assign p31_S0__203_comb = p30_a__35[1:0] ^ p30_a__35[12:11] ^ p30_a__35[21:20];
  assign p31_S0__202_comb = p30_a__35[31:21] ^ p30_a__35[10:0] ^ p30_a__35[19:9];
  assign p31_S0__201_comb = p30_a__35[20:12] ^ p30_a__35[31:23] ^ p30_a__35[8:0];
  assign p31_S0__200_comb = p30_a__35[11:2] ^ p30_a__35[22:13] ^ p30_a__35[31:22];
  assign p31_and_60701_comb = p30_a__35 & p30_a__34;
  assign p31_s_1__147_comb = p31_value__69_comb[16:7] ^ p31_value__69_comb[18:9];
  assign p31_s_1__146_comb = p31_value__69_comb[6:0] ^ p31_value__69_comb[8:2] ^ p31_value__69_comb[31:25];
  assign p31_s_1__145_comb = p31_value__69_comb[31:30] ^ p31_value__69_comb[1:0] ^ p31_value__69_comb[24:23];
  assign p31_s_1__144_comb = p31_value__69_comb[29:17] ^ p31_value__69_comb[31:19] ^ p31_value__69_comb[22:10];
  assign p31_s_1__167_comb = p30_value__84[16:7] ^ p30_value__84[18:9];
  assign p31_s_1__166_comb = p30_value__84[6:0] ^ p30_value__84[8:2] ^ p30_value__84[31:25];
  assign p31_s_1__165_comb = p30_value__84[31:30] ^ p30_value__84[1:0] ^ p30_value__84[24:23];
  assign p31_s_1__164_comb = p30_value__84[29:17] ^ p30_value__84[31:19] ^ p30_value__84[22:10];
  assign p31_S1__207_comb = p31_e__36_comb[5:0] ^ p31_e__36_comb[10:5] ^ p31_e__36_comb[24:19];
  assign p31_S1__206_comb = p31_e__36_comb[31:27] ^ p31_e__36_comb[4:0] ^ p31_e__36_comb[18:14];
  assign p31_S1__205_comb = p31_e__36_comb[26:13] ^ p31_e__36_comb[31:18] ^ p31_e__36_comb[13:0];
  assign p31_S1__204_comb = p31_e__36_comb[12:6] ^ p31_e__36_comb[17:11] ^ p31_e__36_comb[31:25];
  assign p31_add_60661_comb = p30_value__63[31:2] + 30'h1942_9cd5;
  assign p31_S0__35_comb = {p31_S0__203_comb, p31_S0__202_comb, p31_S0__201_comb, p31_S0__200_comb};
  assign p31_maj__35_comb = p31_and_60701_comb ^ p30_a__35 & p30_a__33 ^ p30_and_60523;
  assign p31_s_1__25_comb = {p31_s_1__147_comb, p31_s_1__146_comb, p31_s_1__145_comb, p31_s_1__144_comb};
  assign p31_s_1__30_comb = {p31_s_1__167_comb, p31_s_1__166_comb, p31_s_1__165_comb, p31_s_1__164_comb};
  assign p31_s_0__175_comb = p30_value__51[6:4] ^ p30_value__51[17:15];
  assign p31_s_0__174_comb = p30_value__51[3:0] ^ p30_value__51[14:11] ^ p30_value__51[31:28];
  assign p31_s_0__173_comb = p30_value__51[31:21] ^ p30_value__51[10:0] ^ p30_value__51[27:17];
  assign p31_s_0__172_comb = p30_value__51[20:7] ^ p30_value__51[31:18] ^ p30_value__51[16:3];
  assign p31_s_0__179_comb = p30_value__54[6:4] ^ p30_value__54[17:15];
  assign p31_s_0__178_comb = p30_value__54[3:0] ^ p30_value__54[14:11] ^ p30_value__54[31:28];
  assign p31_s_0__177_comb = p30_value__54[31:21] ^ p30_value__54[10:0] ^ p30_value__54[27:17];
  assign p31_s_0__176_comb = p30_value__54[20:7] ^ p30_value__54[31:18] ^ p30_value__54[16:3];
  assign p31_s_0__183_comb = p30_value__57[6:4] ^ p30_value__57[17:15];
  assign p31_s_0__182_comb = p30_value__57[3:0] ^ p30_value__57[14:11] ^ p30_value__57[31:28];
  assign p31_s_0__181_comb = p30_value__57[31:21] ^ p30_value__57[10:0] ^ p30_value__57[27:17];
  assign p31_s_0__180_comb = p30_value__57[20:7] ^ p30_value__57[31:18] ^ p30_value__57[16:3];
  assign p31_s_0__187_comb = p30_value__60[6:4] ^ p30_value__60[17:15];
  assign p31_s_0__186_comb = p30_value__60[3:0] ^ p30_value__60[14:11] ^ p30_value__60[31:28];
  assign p31_s_0__185_comb = p30_value__60[31:21] ^ p30_value__60[10:0] ^ p30_value__60[27:17];
  assign p31_s_0__184_comb = p30_value__60[20:7] ^ p30_value__60[31:18] ^ p30_value__60[16:3];
  assign p31_S1__36_comb = {p31_S1__207_comb, p31_S1__206_comb, p31_S1__205_comb, p31_S1__204_comb};
  assign p31_ch__36_comb = p31_e__36_comb & p30_e__35 ^ ~(p31_e__36_comb | ~p30_e__34);
  assign p31_temp1__294_comb = {p31_add_60661_comb, p30_value__63[1:0]};
  assign p31_temp2__35_comb = p31_S0__35_comb + p31_maj__35_comb;
  assign p31_value__74_comb = p30_value__54 + p31_s_1__25_comb;
  assign p31_value__89_comb = p31_value__69_comb + p31_s_1__30_comb;
  assign p31_s_0__32_comb = {p31_s_0__175_comb, p31_s_0__174_comb, p31_s_0__173_comb, p31_s_0__172_comb};
  assign p31_s_0__33_comb = {p31_s_0__179_comb, p31_s_0__178_comb, p31_s_0__177_comb, p31_s_0__176_comb};
  assign p31_s_0__34_comb = {p31_s_0__183_comb, p31_s_0__182_comb, p31_s_0__181_comb, p31_s_0__180_comb};
  assign p31_s_0__35_comb = {p31_s_0__187_comb, p31_s_0__186_comb, p31_s_0__185_comb, p31_s_0__184_comb};
  assign p31_temp1__389_comb = p30_e__33 + p31_S1__36_comb;
  assign p31_temp1__390_comb = p31_ch__36_comb + p31_temp1__294_comb;
  assign p31_a__36_comb = p31_temp1__144_comb + p31_temp2__35_comb;
  assign p31_value__75_comb = p30_value__73 + p31_value__74_comb;
  assign p31_value__90_comb = p30_value__88 + p31_value__89_comb;
  assign p31_value__94_comb = p30_value__48 + p31_s_0__32_comb;
  assign p31_value__97_comb = p30_value__51 + p31_s_0__33_comb;
  assign p31_value__100_comb = p30_value__54 + p31_s_0__34_comb;
  assign p31_value__103_comb = p30_value__57 + p31_s_0__35_comb;

  // Registers for pipe stage 31:
  reg [31:0] p31_e__34;
  reg [31:0] p31_e__35;
  reg [31:0] p31_value__60;
  reg [31:0] p31_e__36;
  reg [31:0] p31_value__63;
  reg [31:0] p31_temp1__389;
  reg [31:0] p31_temp1__390;
  reg [31:0] p31_a__33;
  reg [31:0] p31_value__66;
  reg [31:0] p31_a__34;
  reg [31:0] p31_value__69;
  reg [31:0] p31_a__35;
  reg [31:0] p31_and_60701;
  reg [31:0] p31_value__72;
  reg [31:0] p31_a__36;
  reg [31:0] p31_value__75;
  reg [31:0] p31_value__78;
  reg [31:0] p31_value__79;
  reg [31:0] p31_value__84;
  reg [31:0] p31_value__85;
  reg [31:0] p31_value__90;
  reg [31:0] p31_value__91;
  reg [31:0] p31_value__94;
  reg [31:0] p31_value__97;
  reg [31:0] p31_value__100;
  reg [31:0] p31_value__103;
  always_ff @ (posedge clk) begin
    p31_e__34 <= p30_e__34;
    p31_e__35 <= p30_e__35;
    p31_value__60 <= p30_value__60;
    p31_e__36 <= p31_e__36_comb;
    p31_value__63 <= p30_value__63;
    p31_temp1__389 <= p31_temp1__389_comb;
    p31_temp1__390 <= p31_temp1__390_comb;
    p31_a__33 <= p30_a__33;
    p31_value__66 <= p30_value__66;
    p31_a__34 <= p30_a__34;
    p31_value__69 <= p31_value__69_comb;
    p31_a__35 <= p30_a__35;
    p31_and_60701 <= p31_and_60701_comb;
    p31_value__72 <= p30_value__72;
    p31_a__36 <= p31_a__36_comb;
    p31_value__75 <= p31_value__75_comb;
    p31_value__78 <= p30_value__78;
    p31_value__79 <= p30_value__79;
    p31_value__84 <= p30_value__84;
    p31_value__85 <= p30_value__85;
    p31_value__90 <= p31_value__90_comb;
    p31_value__91 <= p30_value__91;
    p31_value__94 <= p31_value__94_comb;
    p31_value__97 <= p31_value__97_comb;
    p31_value__100 <= p31_value__100_comb;
    p31_value__103 <= p31_value__103_comb;
  end

  // ===== Pipe stage 32:
  wire [9:0] p32_s_1__155_comb;
  wire [6:0] p32_s_1__154_comb;
  wire [1:0] p32_s_1__153_comb;
  wire [12:0] p32_s_1__152_comb;
  wire [31:0] p32_s_1__27_comb;
  wire [31:0] p32_temp1__391_comb;
  wire [31:0] p32_value__80_comb;
  wire [31:0] p32_e__37_comb;
  wire [31:0] p32_value__81_comb;
  wire [5:0] p32_S1__211_comb;
  wire [4:0] p32_S1__210_comb;
  wire [13:0] p32_S1__209_comb;
  wire [6:0] p32_S1__208_comb;
  wire [1:0] p32_S0__207_comb;
  wire [10:0] p32_S0__206_comb;
  wire [8:0] p32_S0__205_comb;
  wire [9:0] p32_S0__204_comb;
  wire [31:0] p32_and_60906_comb;
  wire [9:0] p32_s_1__163_comb;
  wire [6:0] p32_s_1__162_comb;
  wire [1:0] p32_s_1__161_comb;
  wire [12:0] p32_s_1__160_comb;
  wire [31:0] p32_S1__37_comb;
  wire [31:0] p32_S0__36_comb;
  wire [31:0] p32_maj__36_comb;
  wire [31:0] p32_s_1__29_comb;
  wire [2:0] p32_s_0__191_comb;
  wire [3:0] p32_s_0__190_comb;
  wire [10:0] p32_s_0__189_comb;
  wire [13:0] p32_s_0__188_comb;
  wire [2:0] p32_s_0__195_comb;
  wire [3:0] p32_s_0__194_comb;
  wire [10:0] p32_s_0__193_comb;
  wire [13:0] p32_s_0__192_comb;
  wire [2:0] p32_s_0__199_comb;
  wire [3:0] p32_s_0__198_comb;
  wire [10:0] p32_s_0__197_comb;
  wire [13:0] p32_s_0__196_comb;
  wire [31:0] p32_temp1__149_comb;
  wire [31:0] p32_ch__37_comb;
  wire [31:0] p32_temp2__36_comb;
  wire [31:0] p32_value__86_comb;
  wire [31:0] p32_s_0__36_comb;
  wire [31:0] p32_s_0__37_comb;
  wire [31:0] p32_s_0__38_comb;
  wire [31:0] p32_temp1__150_comb;
  wire [31:0] p32_temp1__295_comb;
  wire [31:0] p32_a__37_comb;
  wire [31:0] p32_value__87_comb;
  wire [31:0] p32_value__106_comb;
  wire [31:0] p32_value__109_comb;
  wire [31:0] p32_value__112_comb;
  assign p32_s_1__155_comb = p31_value__75[16:7] ^ p31_value__75[18:9];
  assign p32_s_1__154_comb = p31_value__75[6:0] ^ p31_value__75[8:2] ^ p31_value__75[31:25];
  assign p32_s_1__153_comb = p31_value__75[31:30] ^ p31_value__75[1:0] ^ p31_value__75[24:23];
  assign p32_s_1__152_comb = p31_value__75[29:17] ^ p31_value__75[31:19] ^ p31_value__75[22:10];
  assign p32_s_1__27_comb = {p32_s_1__155_comb, p32_s_1__154_comb, p32_s_1__153_comb, p32_s_1__152_comb};
  assign p32_temp1__391_comb = p31_temp1__389 + p31_temp1__390;
  assign p32_value__80_comb = p31_value__60 + p32_s_1__27_comb;
  assign p32_e__37_comb = p31_a__33 + p32_temp1__391_comb;
  assign p32_value__81_comb = p31_value__79 + p32_value__80_comb;
  assign p32_S1__211_comb = p32_e__37_comb[5:0] ^ p32_e__37_comb[10:5] ^ p32_e__37_comb[24:19];
  assign p32_S1__210_comb = p32_e__37_comb[31:27] ^ p32_e__37_comb[4:0] ^ p32_e__37_comb[18:14];
  assign p32_S1__209_comb = p32_e__37_comb[26:13] ^ p32_e__37_comb[31:18] ^ p32_e__37_comb[13:0];
  assign p32_S1__208_comb = p32_e__37_comb[12:6] ^ p32_e__37_comb[17:11] ^ p32_e__37_comb[31:25];
  assign p32_S0__207_comb = p31_a__36[1:0] ^ p31_a__36[12:11] ^ p31_a__36[21:20];
  assign p32_S0__206_comb = p31_a__36[31:21] ^ p31_a__36[10:0] ^ p31_a__36[19:9];
  assign p32_S0__205_comb = p31_a__36[20:12] ^ p31_a__36[31:23] ^ p31_a__36[8:0];
  assign p32_S0__204_comb = p31_a__36[11:2] ^ p31_a__36[22:13] ^ p31_a__36[31:22];
  assign p32_and_60906_comb = p31_a__36 & p31_a__35;
  assign p32_s_1__163_comb = p32_value__81_comb[16:7] ^ p32_value__81_comb[18:9];
  assign p32_s_1__162_comb = p32_value__81_comb[6:0] ^ p32_value__81_comb[8:2] ^ p32_value__81_comb[31:25];
  assign p32_s_1__161_comb = p32_value__81_comb[31:30] ^ p32_value__81_comb[1:0] ^ p32_value__81_comb[24:23];
  assign p32_s_1__160_comb = p32_value__81_comb[29:17] ^ p32_value__81_comb[31:19] ^ p32_value__81_comb[22:10];
  assign p32_S1__37_comb = {p32_S1__211_comb, p32_S1__210_comb, p32_S1__209_comb, p32_S1__208_comb};
  assign p32_S0__36_comb = {p32_S0__207_comb, p32_S0__206_comb, p32_S0__205_comb, p32_S0__204_comb};
  assign p32_maj__36_comb = p32_and_60906_comb ^ p31_a__36 & p31_a__34 ^ p31_and_60701;
  assign p32_s_1__29_comb = {p32_s_1__163_comb, p32_s_1__162_comb, p32_s_1__161_comb, p32_s_1__160_comb};
  assign p32_s_0__191_comb = p31_value__63[6:4] ^ p31_value__63[17:15];
  assign p32_s_0__190_comb = p31_value__63[3:0] ^ p31_value__63[14:11] ^ p31_value__63[31:28];
  assign p32_s_0__189_comb = p31_value__63[31:21] ^ p31_value__63[10:0] ^ p31_value__63[27:17];
  assign p32_s_0__188_comb = p31_value__63[20:7] ^ p31_value__63[31:18] ^ p31_value__63[16:3];
  assign p32_s_0__195_comb = p31_value__66[6:4] ^ p31_value__66[17:15];
  assign p32_s_0__194_comb = p31_value__66[3:0] ^ p31_value__66[14:11] ^ p31_value__66[31:28];
  assign p32_s_0__193_comb = p31_value__66[31:21] ^ p31_value__66[10:0] ^ p31_value__66[27:17];
  assign p32_s_0__192_comb = p31_value__66[20:7] ^ p31_value__66[31:18] ^ p31_value__66[16:3];
  assign p32_s_0__199_comb = p31_value__69[6:4] ^ p31_value__69[17:15];
  assign p32_s_0__198_comb = p31_value__69[3:0] ^ p31_value__69[14:11] ^ p31_value__69[31:28];
  assign p32_s_0__197_comb = p31_value__69[31:21] ^ p31_value__69[10:0] ^ p31_value__69[27:17];
  assign p32_s_0__196_comb = p31_value__69[20:7] ^ p31_value__69[31:18] ^ p31_value__69[16:3];
  assign p32_temp1__149_comb = p31_e__34 + p32_S1__37_comb;
  assign p32_ch__37_comb = p32_e__37_comb & p31_e__36 ^ ~(p32_e__37_comb | ~p31_e__35);
  assign p32_temp2__36_comb = p32_S0__36_comb + p32_maj__36_comb;
  assign p32_value__86_comb = p31_value__66 + p32_s_1__29_comb;
  assign p32_s_0__36_comb = {p32_s_0__191_comb, p32_s_0__190_comb, p32_s_0__189_comb, p32_s_0__188_comb};
  assign p32_s_0__37_comb = {p32_s_0__195_comb, p32_s_0__194_comb, p32_s_0__193_comb, p32_s_0__192_comb};
  assign p32_s_0__38_comb = {p32_s_0__199_comb, p32_s_0__198_comb, p32_s_0__197_comb, p32_s_0__196_comb};
  assign p32_temp1__150_comb = p32_temp1__149_comb + p32_ch__37_comb;
  assign p32_temp1__295_comb = p31_value__66 + 32'h766a_0abb;
  assign p32_a__37_comb = p32_temp1__391_comb + p32_temp2__36_comb;
  assign p32_value__87_comb = p31_value__85 + p32_value__86_comb;
  assign p32_value__106_comb = p31_value__60 + p32_s_0__36_comb;
  assign p32_value__109_comb = p31_value__63 + p32_s_0__37_comb;
  assign p32_value__112_comb = p31_value__66 + p32_s_0__38_comb;

  // Registers for pipe stage 32:
  reg [31:0] p32_e__35;
  reg [31:0] p32_e__36;
  reg [31:0] p32_e__37;
  reg [31:0] p32_temp1__150;
  reg [31:0] p32_temp1__295;
  reg [31:0] p32_a__34;
  reg [31:0] p32_value__69;
  reg [31:0] p32_a__35;
  reg [31:0] p32_value__72;
  reg [31:0] p32_a__36;
  reg [31:0] p32_and_60906;
  reg [31:0] p32_value__75;
  reg [31:0] p32_a__37;
  reg [31:0] p32_value__78;
  reg [31:0] p32_value__81;
  reg [31:0] p32_value__84;
  reg [31:0] p32_value__87;
  reg [31:0] p32_value__90;
  reg [31:0] p32_value__91;
  reg [31:0] p32_value__94;
  reg [31:0] p32_value__97;
  reg [31:0] p32_value__100;
  reg [31:0] p32_value__103;
  reg [31:0] p32_value__106;
  reg [31:0] p32_value__109;
  reg [31:0] p32_value__112;
  always_ff @ (posedge clk) begin
    p32_e__35 <= p31_e__35;
    p32_e__36 <= p31_e__36;
    p32_e__37 <= p32_e__37_comb;
    p32_temp1__150 <= p32_temp1__150_comb;
    p32_temp1__295 <= p32_temp1__295_comb;
    p32_a__34 <= p31_a__34;
    p32_value__69 <= p31_value__69;
    p32_a__35 <= p31_a__35;
    p32_value__72 <= p31_value__72;
    p32_a__36 <= p31_a__36;
    p32_and_60906 <= p32_and_60906_comb;
    p32_value__75 <= p31_value__75;
    p32_a__37 <= p32_a__37_comb;
    p32_value__78 <= p31_value__78;
    p32_value__81 <= p32_value__81_comb;
    p32_value__84 <= p31_value__84;
    p32_value__87 <= p32_value__87_comb;
    p32_value__90 <= p31_value__90;
    p32_value__91 <= p31_value__91;
    p32_value__94 <= p31_value__94;
    p32_value__97 <= p31_value__97;
    p32_value__100 <= p31_value__100;
    p32_value__103 <= p31_value__103;
    p32_value__106 <= p32_value__106_comb;
    p32_value__109 <= p32_value__109_comb;
    p32_value__112 <= p32_value__112_comb;
  end

  // ===== Pipe stage 33:
  wire [9:0] p33_s_1__171_comb;
  wire [6:0] p33_s_1__170_comb;
  wire [1:0] p33_s_1__169_comb;
  wire [12:0] p33_s_1__168_comb;
  wire [31:0] p33_s_1__31_comb;
  wire [31:0] p33_temp1__152_comb;
  wire [31:0] p33_value__92_comb;
  wire [31:0] p33_e__38_comb;
  wire [31:0] p33_value__93_comb;
  wire [5:0] p33_S1__215_comb;
  wire [4:0] p33_S1__214_comb;
  wire [13:0] p33_S1__213_comb;
  wire [6:0] p33_S1__212_comb;
  wire [30:0] p33_add_61074_comb;
  wire [1:0] p33_S0__211_comb;
  wire [10:0] p33_S0__210_comb;
  wire [8:0] p33_S0__209_comb;
  wire [9:0] p33_S0__208_comb;
  wire [31:0] p33_and_61098_comb;
  wire [9:0] p33_s_1__179_comb;
  wire [6:0] p33_s_1__178_comb;
  wire [1:0] p33_s_1__177_comb;
  wire [12:0] p33_s_1__176_comb;
  wire [31:0] p33_S1__38_comb;
  wire [31:0] p33_ch__38_comb;
  wire [31:0] p33_temp1__296_comb;
  wire [31:0] p33_S0__37_comb;
  wire [31:0] p33_maj__37_comb;
  wire [31:0] p33_s_1__33_comb;
  wire [2:0] p33_s_0__203_comb;
  wire [3:0] p33_s_0__202_comb;
  wire [10:0] p33_s_0__201_comb;
  wire [13:0] p33_s_0__200_comb;
  wire [31:0] p33_temp1__386_comb;
  wire [31:0] p33_temp1__387_comb;
  wire [31:0] p33_temp2__37_comb;
  wire [31:0] p33_value__98_comb;
  wire [31:0] p33_s_0__39_comb;
  wire [31:0] p33_temp1__388_comb;
  wire [31:0] p33_a__38_comb;
  wire [31:0] p33_value__99_comb;
  wire [31:0] p33_value__115_comb;
  assign p33_s_1__171_comb = p32_value__87[16:7] ^ p32_value__87[18:9];
  assign p33_s_1__170_comb = p32_value__87[6:0] ^ p32_value__87[8:2] ^ p32_value__87[31:25];
  assign p33_s_1__169_comb = p32_value__87[31:30] ^ p32_value__87[1:0] ^ p32_value__87[24:23];
  assign p33_s_1__168_comb = p32_value__87[29:17] ^ p32_value__87[31:19] ^ p32_value__87[22:10];
  assign p33_s_1__31_comb = {p33_s_1__171_comb, p33_s_1__170_comb, p33_s_1__169_comb, p33_s_1__168_comb};
  assign p33_temp1__152_comb = p32_temp1__150 + p32_temp1__295;
  assign p33_value__92_comb = p32_value__72 + p33_s_1__31_comb;
  assign p33_e__38_comb = p32_a__34 + p33_temp1__152_comb;
  assign p33_value__93_comb = p32_value__91 + p33_value__92_comb;
  assign p33_S1__215_comb = p33_e__38_comb[5:0] ^ p33_e__38_comb[10:5] ^ p33_e__38_comb[24:19];
  assign p33_S1__214_comb = p33_e__38_comb[31:27] ^ p33_e__38_comb[4:0] ^ p33_e__38_comb[18:14];
  assign p33_S1__213_comb = p33_e__38_comb[26:13] ^ p33_e__38_comb[31:18] ^ p33_e__38_comb[13:0];
  assign p33_S1__212_comb = p33_e__38_comb[12:6] ^ p33_e__38_comb[17:11] ^ p33_e__38_comb[31:25];
  assign p33_add_61074_comb = p32_value__69[31:1] + 31'h40e1_6497;
  assign p33_S0__211_comb = p32_a__37[1:0] ^ p32_a__37[12:11] ^ p32_a__37[21:20];
  assign p33_S0__210_comb = p32_a__37[31:21] ^ p32_a__37[10:0] ^ p32_a__37[19:9];
  assign p33_S0__209_comb = p32_a__37[20:12] ^ p32_a__37[31:23] ^ p32_a__37[8:0];
  assign p33_S0__208_comb = p32_a__37[11:2] ^ p32_a__37[22:13] ^ p32_a__37[31:22];
  assign p33_and_61098_comb = p32_a__37 & p32_a__36;
  assign p33_s_1__179_comb = p33_value__93_comb[16:7] ^ p33_value__93_comb[18:9];
  assign p33_s_1__178_comb = p33_value__93_comb[6:0] ^ p33_value__93_comb[8:2] ^ p33_value__93_comb[31:25];
  assign p33_s_1__177_comb = p33_value__93_comb[31:30] ^ p33_value__93_comb[1:0] ^ p33_value__93_comb[24:23];
  assign p33_s_1__176_comb = p33_value__93_comb[29:17] ^ p33_value__93_comb[31:19] ^ p33_value__93_comb[22:10];
  assign p33_S1__38_comb = {p33_S1__215_comb, p33_S1__214_comb, p33_S1__213_comb, p33_S1__212_comb};
  assign p33_ch__38_comb = p33_e__38_comb & p32_e__37 ^ ~(p33_e__38_comb | ~p32_e__36);
  assign p33_temp1__296_comb = {p33_add_61074_comb, p32_value__69[0]};
  assign p33_S0__37_comb = {p33_S0__211_comb, p33_S0__210_comb, p33_S0__209_comb, p33_S0__208_comb};
  assign p33_maj__37_comb = p33_and_61098_comb ^ p32_a__37 & p32_a__35 ^ p32_and_60906;
  assign p33_s_1__33_comb = {p33_s_1__179_comb, p33_s_1__178_comb, p33_s_1__177_comb, p33_s_1__176_comb};
  assign p33_s_0__203_comb = p32_value__72[6:4] ^ p32_value__72[17:15];
  assign p33_s_0__202_comb = p32_value__72[3:0] ^ p32_value__72[14:11] ^ p32_value__72[31:28];
  assign p33_s_0__201_comb = p32_value__72[31:21] ^ p32_value__72[10:0] ^ p32_value__72[27:17];
  assign p33_s_0__200_comb = p32_value__72[20:7] ^ p32_value__72[31:18] ^ p32_value__72[16:3];
  assign p33_temp1__386_comb = p32_e__35 + p33_S1__38_comb;
  assign p33_temp1__387_comb = p33_ch__38_comb + p33_temp1__296_comb;
  assign p33_temp2__37_comb = p33_S0__37_comb + p33_maj__37_comb;
  assign p33_value__98_comb = p32_value__78 + p33_s_1__33_comb;
  assign p33_s_0__39_comb = {p33_s_0__203_comb, p33_s_0__202_comb, p33_s_0__201_comb, p33_s_0__200_comb};
  assign p33_temp1__388_comb = p33_temp1__386_comb + p33_temp1__387_comb;
  assign p33_a__38_comb = p33_temp1__152_comb + p33_temp2__37_comb;
  assign p33_value__99_comb = p32_value__97 + p33_value__98_comb;
  assign p33_value__115_comb = p32_value__69 + p33_s_0__39_comb;

  // Registers for pipe stage 33:
  reg [31:0] p33_e__36;
  reg [31:0] p33_e__37;
  reg [31:0] p33_e__38;
  reg [31:0] p33_a__35;
  reg [31:0] p33_temp1__388;
  reg [31:0] p33_value__72;
  reg [31:0] p33_a__36;
  reg [31:0] p33_value__75;
  reg [31:0] p33_a__37;
  reg [31:0] p33_and_61098;
  reg [31:0] p33_value__78;
  reg [31:0] p33_a__38;
  reg [31:0] p33_value__81;
  reg [31:0] p33_value__84;
  reg [31:0] p33_value__87;
  reg [31:0] p33_value__90;
  reg [31:0] p33_value__93;
  reg [31:0] p33_value__94;
  reg [31:0] p33_value__99;
  reg [31:0] p33_value__100;
  reg [31:0] p33_value__103;
  reg [31:0] p33_value__106;
  reg [31:0] p33_value__109;
  reg [31:0] p33_value__112;
  reg [31:0] p33_value__115;
  always_ff @ (posedge clk) begin
    p33_e__36 <= p32_e__36;
    p33_e__37 <= p32_e__37;
    p33_e__38 <= p33_e__38_comb;
    p33_a__35 <= p32_a__35;
    p33_temp1__388 <= p33_temp1__388_comb;
    p33_value__72 <= p32_value__72;
    p33_a__36 <= p32_a__36;
    p33_value__75 <= p32_value__75;
    p33_a__37 <= p32_a__37;
    p33_and_61098 <= p33_and_61098_comb;
    p33_value__78 <= p32_value__78;
    p33_a__38 <= p33_a__38_comb;
    p33_value__81 <= p32_value__81;
    p33_value__84 <= p32_value__84;
    p33_value__87 <= p32_value__87;
    p33_value__90 <= p32_value__90;
    p33_value__93 <= p33_value__93_comb;
    p33_value__94 <= p32_value__94;
    p33_value__99 <= p33_value__99_comb;
    p33_value__100 <= p32_value__100;
    p33_value__103 <= p32_value__103;
    p33_value__106 <= p32_value__106;
    p33_value__109 <= p32_value__109;
    p33_value__112 <= p32_value__112;
    p33_value__115 <= p33_value__115_comb;
  end

  // ===== Pipe stage 34:
  wire [31:0] p34_e__39_comb;
  wire [5:0] p34_S1__219_comb;
  wire [4:0] p34_S1__218_comb;
  wire [13:0] p34_S1__217_comb;
  wire [6:0] p34_S1__216_comb;
  wire [31:0] p34_S1__39_comb;
  wire [1:0] p34_S0__215_comb;
  wire [10:0] p34_S0__214_comb;
  wire [8:0] p34_S0__213_comb;
  wire [9:0] p34_S0__212_comb;
  wire [31:0] p34_and_61250_comb;
  wire [9:0] p34_s_1__187_comb;
  wire [6:0] p34_s_1__186_comb;
  wire [1:0] p34_s_1__185_comb;
  wire [12:0] p34_s_1__184_comb;
  wire [31:0] p34_temp1__157_comb;
  wire [31:0] p34_ch__39_comb;
  wire [31:0] p34_S0__38_comb;
  wire [31:0] p34_maj__38_comb;
  wire [31:0] p34_s_1__35_comb;
  wire [2:0] p34_s_0__207_comb;
  wire [3:0] p34_s_0__206_comb;
  wire [10:0] p34_s_0__205_comb;
  wire [13:0] p34_s_0__204_comb;
  wire [31:0] p34_temp1__158_comb;
  wire [31:0] p34_temp1__297_comb;
  wire [31:0] p34_temp2__38_comb;
  wire [31:0] p34_value__104_comb;
  wire [31:0] p34_s_0__40_comb;
  wire [31:0] p34_temp1__160_comb;
  wire [31:0] p34_a__39_comb;
  wire [31:0] p34_value__105_comb;
  wire [31:0] p34_value__118_comb;
  assign p34_e__39_comb = p33_a__35 + p33_temp1__388;
  assign p34_S1__219_comb = p34_e__39_comb[5:0] ^ p34_e__39_comb[10:5] ^ p34_e__39_comb[24:19];
  assign p34_S1__218_comb = p34_e__39_comb[31:27] ^ p34_e__39_comb[4:0] ^ p34_e__39_comb[18:14];
  assign p34_S1__217_comb = p34_e__39_comb[26:13] ^ p34_e__39_comb[31:18] ^ p34_e__39_comb[13:0];
  assign p34_S1__216_comb = p34_e__39_comb[12:6] ^ p34_e__39_comb[17:11] ^ p34_e__39_comb[31:25];
  assign p34_S1__39_comb = {p34_S1__219_comb, p34_S1__218_comb, p34_S1__217_comb, p34_S1__216_comb};
  assign p34_S0__215_comb = p33_a__38[1:0] ^ p33_a__38[12:11] ^ p33_a__38[21:20];
  assign p34_S0__214_comb = p33_a__38[31:21] ^ p33_a__38[10:0] ^ p33_a__38[19:9];
  assign p34_S0__213_comb = p33_a__38[20:12] ^ p33_a__38[31:23] ^ p33_a__38[8:0];
  assign p34_S0__212_comb = p33_a__38[11:2] ^ p33_a__38[22:13] ^ p33_a__38[31:22];
  assign p34_and_61250_comb = p33_a__38 & p33_a__37;
  assign p34_s_1__187_comb = p33_value__99[16:7] ^ p33_value__99[18:9];
  assign p34_s_1__186_comb = p33_value__99[6:0] ^ p33_value__99[8:2] ^ p33_value__99[31:25];
  assign p34_s_1__185_comb = p33_value__99[31:30] ^ p33_value__99[1:0] ^ p33_value__99[24:23];
  assign p34_s_1__184_comb = p33_value__99[29:17] ^ p33_value__99[31:19] ^ p33_value__99[22:10];
  assign p34_temp1__157_comb = p33_e__36 + p34_S1__39_comb;
  assign p34_ch__39_comb = p34_e__39_comb & p33_e__38 ^ ~(p34_e__39_comb | ~p33_e__37);
  assign p34_S0__38_comb = {p34_S0__215_comb, p34_S0__214_comb, p34_S0__213_comb, p34_S0__212_comb};
  assign p34_maj__38_comb = p34_and_61250_comb ^ p33_a__38 & p33_a__36 ^ p33_and_61098;
  assign p34_s_1__35_comb = {p34_s_1__187_comb, p34_s_1__186_comb, p34_s_1__185_comb, p34_s_1__184_comb};
  assign p34_s_0__207_comb = p33_value__75[6:4] ^ p33_value__75[17:15];
  assign p34_s_0__206_comb = p33_value__75[3:0] ^ p33_value__75[14:11] ^ p33_value__75[31:28];
  assign p34_s_0__205_comb = p33_value__75[31:21] ^ p33_value__75[10:0] ^ p33_value__75[27:17];
  assign p34_s_0__204_comb = p33_value__75[20:7] ^ p33_value__75[31:18] ^ p33_value__75[16:3];
  assign p34_temp1__158_comb = p34_temp1__157_comb + p34_ch__39_comb;
  assign p34_temp1__297_comb = p33_value__72 + 32'h9272_2c85;
  assign p34_temp2__38_comb = p34_S0__38_comb + p34_maj__38_comb;
  assign p34_value__104_comb = p33_value__84 + p34_s_1__35_comb;
  assign p34_s_0__40_comb = {p34_s_0__207_comb, p34_s_0__206_comb, p34_s_0__205_comb, p34_s_0__204_comb};
  assign p34_temp1__160_comb = p34_temp1__158_comb + p34_temp1__297_comb;
  assign p34_a__39_comb = p33_temp1__388 + p34_temp2__38_comb;
  assign p34_value__105_comb = p33_value__103 + p34_value__104_comb;
  assign p34_value__118_comb = p33_value__72 + p34_s_0__40_comb;

  // Registers for pipe stage 34:
  reg [31:0] p34_e__37;
  reg [31:0] p34_e__38;
  reg [31:0] p34_e__39;
  reg [31:0] p34_a__36;
  reg [31:0] p34_temp1__160;
  reg [31:0] p34_value__75;
  reg [31:0] p34_a__37;
  reg [31:0] p34_value__78;
  reg [31:0] p34_a__38;
  reg [31:0] p34_value__81;
  reg [31:0] p34_and_61250;
  reg [31:0] p34_a__39;
  reg [31:0] p34_value__84;
  reg [31:0] p34_value__87;
  reg [31:0] p34_value__90;
  reg [31:0] p34_value__93;
  reg [31:0] p34_value__94;
  reg [31:0] p34_value__99;
  reg [31:0] p34_value__100;
  reg [31:0] p34_value__105;
  reg [31:0] p34_value__106;
  reg [31:0] p34_value__109;
  reg [31:0] p34_value__112;
  reg [31:0] p34_value__115;
  reg [31:0] p34_value__118;
  always_ff @ (posedge clk) begin
    p34_e__37 <= p33_e__37;
    p34_e__38 <= p33_e__38;
    p34_e__39 <= p34_e__39_comb;
    p34_a__36 <= p33_a__36;
    p34_temp1__160 <= p34_temp1__160_comb;
    p34_value__75 <= p33_value__75;
    p34_a__37 <= p33_a__37;
    p34_value__78 <= p33_value__78;
    p34_a__38 <= p33_a__38;
    p34_value__81 <= p33_value__81;
    p34_and_61250 <= p34_and_61250_comb;
    p34_a__39 <= p34_a__39_comb;
    p34_value__84 <= p33_value__84;
    p34_value__87 <= p33_value__87;
    p34_value__90 <= p33_value__90;
    p34_value__93 <= p33_value__93;
    p34_value__94 <= p33_value__94;
    p34_value__99 <= p33_value__99;
    p34_value__100 <= p33_value__100;
    p34_value__105 <= p34_value__105_comb;
    p34_value__106 <= p33_value__106;
    p34_value__109 <= p33_value__109;
    p34_value__112 <= p33_value__112;
    p34_value__115 <= p33_value__115;
    p34_value__118 <= p34_value__118_comb;
  end

  // ===== Pipe stage 35:
  wire [31:0] p35_e__40_comb;
  wire [5:0] p35_S1__223_comb;
  wire [4:0] p35_S1__222_comb;
  wire [13:0] p35_S1__221_comb;
  wire [6:0] p35_S1__220_comb;
  wire [31:0] p35_S1__40_comb;
  wire [1:0] p35_S0__219_comb;
  wire [10:0] p35_S0__218_comb;
  wire [8:0] p35_S0__217_comb;
  wire [9:0] p35_S0__216_comb;
  wire [31:0] p35_and_61384_comb;
  wire [31:0] p35_temp1__161_comb;
  wire [31:0] p35_ch__40_comb;
  wire [31:0] p35_S0__39_comb;
  wire [31:0] p35_maj__39_comb;
  wire [31:0] p35_temp1__162_comb;
  wire [31:0] p35_temp1__298_comb;
  wire [31:0] p35_temp2__39_comb;
  wire [31:0] p35_temp1__164_comb;
  wire [31:0] p35_a__40_comb;
  assign p35_e__40_comb = p34_a__36 + p34_temp1__160;
  assign p35_S1__223_comb = p35_e__40_comb[5:0] ^ p35_e__40_comb[10:5] ^ p35_e__40_comb[24:19];
  assign p35_S1__222_comb = p35_e__40_comb[31:27] ^ p35_e__40_comb[4:0] ^ p35_e__40_comb[18:14];
  assign p35_S1__221_comb = p35_e__40_comb[26:13] ^ p35_e__40_comb[31:18] ^ p35_e__40_comb[13:0];
  assign p35_S1__220_comb = p35_e__40_comb[12:6] ^ p35_e__40_comb[17:11] ^ p35_e__40_comb[31:25];
  assign p35_S1__40_comb = {p35_S1__223_comb, p35_S1__222_comb, p35_S1__221_comb, p35_S1__220_comb};
  assign p35_S0__219_comb = p34_a__39[1:0] ^ p34_a__39[12:11] ^ p34_a__39[21:20];
  assign p35_S0__218_comb = p34_a__39[31:21] ^ p34_a__39[10:0] ^ p34_a__39[19:9];
  assign p35_S0__217_comb = p34_a__39[20:12] ^ p34_a__39[31:23] ^ p34_a__39[8:0];
  assign p35_S0__216_comb = p34_a__39[11:2] ^ p34_a__39[22:13] ^ p34_a__39[31:22];
  assign p35_and_61384_comb = p34_a__39 & p34_a__38;
  assign p35_temp1__161_comb = p34_e__37 + p35_S1__40_comb;
  assign p35_ch__40_comb = p35_e__40_comb & p34_e__39 ^ ~(p35_e__40_comb | ~p34_e__38);
  assign p35_S0__39_comb = {p35_S0__219_comb, p35_S0__218_comb, p35_S0__217_comb, p35_S0__216_comb};
  assign p35_maj__39_comb = p35_and_61384_comb ^ p34_a__39 & p34_a__37 ^ p34_and_61250;
  assign p35_temp1__162_comb = p35_temp1__161_comb + p35_ch__40_comb;
  assign p35_temp1__298_comb = p34_value__75 + 32'ha2bf_e8a1;
  assign p35_temp2__39_comb = p35_S0__39_comb + p35_maj__39_comb;
  assign p35_temp1__164_comb = p35_temp1__162_comb + p35_temp1__298_comb;
  assign p35_a__40_comb = p34_temp1__160 + p35_temp2__39_comb;

  // Registers for pipe stage 35:
  reg [31:0] p35_e__38;
  reg [31:0] p35_e__39;
  reg [31:0] p35_e__40;
  reg [31:0] p35_value__75;
  reg [31:0] p35_a__37;
  reg [31:0] p35_temp1__164;
  reg [31:0] p35_value__78;
  reg [31:0] p35_a__38;
  reg [31:0] p35_value__81;
  reg [31:0] p35_a__39;
  reg [31:0] p35_and_61384;
  reg [31:0] p35_value__84;
  reg [31:0] p35_a__40;
  reg [31:0] p35_value__87;
  reg [31:0] p35_value__90;
  reg [31:0] p35_value__93;
  reg [31:0] p35_value__94;
  reg [31:0] p35_value__99;
  reg [31:0] p35_value__100;
  reg [31:0] p35_value__105;
  reg [31:0] p35_value__106;
  reg [31:0] p35_value__109;
  reg [31:0] p35_value__112;
  reg [31:0] p35_value__115;
  reg [31:0] p35_value__118;
  always_ff @ (posedge clk) begin
    p35_e__38 <= p34_e__38;
    p35_e__39 <= p34_e__39;
    p35_e__40 <= p35_e__40_comb;
    p35_value__75 <= p34_value__75;
    p35_a__37 <= p34_a__37;
    p35_temp1__164 <= p35_temp1__164_comb;
    p35_value__78 <= p34_value__78;
    p35_a__38 <= p34_a__38;
    p35_value__81 <= p34_value__81;
    p35_a__39 <= p34_a__39;
    p35_and_61384 <= p35_and_61384_comb;
    p35_value__84 <= p34_value__84;
    p35_a__40 <= p35_a__40_comb;
    p35_value__87 <= p34_value__87;
    p35_value__90 <= p34_value__90;
    p35_value__93 <= p34_value__93;
    p35_value__94 <= p34_value__94;
    p35_value__99 <= p34_value__99;
    p35_value__100 <= p34_value__100;
    p35_value__105 <= p34_value__105;
    p35_value__106 <= p34_value__106;
    p35_value__109 <= p34_value__109;
    p35_value__112 <= p34_value__112;
    p35_value__115 <= p34_value__115;
    p35_value__118 <= p34_value__118;
  end

  // ===== Pipe stage 36:
  wire [31:0] p36_e__41_comb;
  wire [5:0] p36_S1__227_comb;
  wire [4:0] p36_S1__226_comb;
  wire [13:0] p36_S1__225_comb;
  wire [6:0] p36_S1__224_comb;
  wire [31:0] p36_S1__41_comb;
  wire [1:0] p36_S0__223_comb;
  wire [10:0] p36_S0__222_comb;
  wire [8:0] p36_S0__221_comb;
  wire [9:0] p36_S0__220_comb;
  wire [31:0] p36_and_61483_comb;
  wire [31:0] p36_temp1__165_comb;
  wire [31:0] p36_ch__41_comb;
  wire [31:0] p36_S0__40_comb;
  wire [31:0] p36_maj__40_comb;
  wire [31:0] p36_temp1__166_comb;
  wire [31:0] p36_temp1__299_comb;
  wire [31:0] p36_temp2__40_comb;
  wire [31:0] p36_temp1__168_comb;
  wire [31:0] p36_a__41_comb;
  assign p36_e__41_comb = p35_a__37 + p35_temp1__164;
  assign p36_S1__227_comb = p36_e__41_comb[5:0] ^ p36_e__41_comb[10:5] ^ p36_e__41_comb[24:19];
  assign p36_S1__226_comb = p36_e__41_comb[31:27] ^ p36_e__41_comb[4:0] ^ p36_e__41_comb[18:14];
  assign p36_S1__225_comb = p36_e__41_comb[26:13] ^ p36_e__41_comb[31:18] ^ p36_e__41_comb[13:0];
  assign p36_S1__224_comb = p36_e__41_comb[12:6] ^ p36_e__41_comb[17:11] ^ p36_e__41_comb[31:25];
  assign p36_S1__41_comb = {p36_S1__227_comb, p36_S1__226_comb, p36_S1__225_comb, p36_S1__224_comb};
  assign p36_S0__223_comb = p35_a__40[1:0] ^ p35_a__40[12:11] ^ p35_a__40[21:20];
  assign p36_S0__222_comb = p35_a__40[31:21] ^ p35_a__40[10:0] ^ p35_a__40[19:9];
  assign p36_S0__221_comb = p35_a__40[20:12] ^ p35_a__40[31:23] ^ p35_a__40[8:0];
  assign p36_S0__220_comb = p35_a__40[11:2] ^ p35_a__40[22:13] ^ p35_a__40[31:22];
  assign p36_and_61483_comb = p35_a__40 & p35_a__39;
  assign p36_temp1__165_comb = p35_e__38 + p36_S1__41_comb;
  assign p36_ch__41_comb = p36_e__41_comb & p35_e__40 ^ ~(p36_e__41_comb | ~p35_e__39);
  assign p36_S0__40_comb = {p36_S0__223_comb, p36_S0__222_comb, p36_S0__221_comb, p36_S0__220_comb};
  assign p36_maj__40_comb = p36_and_61483_comb ^ p35_a__40 & p35_a__38 ^ p35_and_61384;
  assign p36_temp1__166_comb = p36_temp1__165_comb + p36_ch__41_comb;
  assign p36_temp1__299_comb = p35_value__78 + 32'ha81a_664b;
  assign p36_temp2__40_comb = p36_S0__40_comb + p36_maj__40_comb;
  assign p36_temp1__168_comb = p36_temp1__166_comb + p36_temp1__299_comb;
  assign p36_a__41_comb = p35_temp1__164 + p36_temp2__40_comb;

  // Registers for pipe stage 36:
  reg [31:0] p36_e__39;
  reg [31:0] p36_e__40;
  reg [31:0] p36_value__75;
  reg [31:0] p36_e__41;
  reg [31:0] p36_value__78;
  reg [31:0] p36_a__38;
  reg [31:0] p36_temp1__168;
  reg [31:0] p36_value__81;
  reg [31:0] p36_a__39;
  reg [31:0] p36_value__84;
  reg [31:0] p36_a__40;
  reg [31:0] p36_and_61483;
  reg [31:0] p36_value__87;
  reg [31:0] p36_a__41;
  reg [31:0] p36_value__90;
  reg [31:0] p36_value__93;
  reg [31:0] p36_value__94;
  reg [31:0] p36_value__99;
  reg [31:0] p36_value__100;
  reg [31:0] p36_value__105;
  reg [31:0] p36_value__106;
  reg [31:0] p36_value__109;
  reg [31:0] p36_value__112;
  reg [31:0] p36_value__115;
  reg [31:0] p36_value__118;
  always_ff @ (posedge clk) begin
    p36_e__39 <= p35_e__39;
    p36_e__40 <= p35_e__40;
    p36_value__75 <= p35_value__75;
    p36_e__41 <= p36_e__41_comb;
    p36_value__78 <= p35_value__78;
    p36_a__38 <= p35_a__38;
    p36_temp1__168 <= p36_temp1__168_comb;
    p36_value__81 <= p35_value__81;
    p36_a__39 <= p35_a__39;
    p36_value__84 <= p35_value__84;
    p36_a__40 <= p35_a__40;
    p36_and_61483 <= p36_and_61483_comb;
    p36_value__87 <= p35_value__87;
    p36_a__41 <= p36_a__41_comb;
    p36_value__90 <= p35_value__90;
    p36_value__93 <= p35_value__93;
    p36_value__94 <= p35_value__94;
    p36_value__99 <= p35_value__99;
    p36_value__100 <= p35_value__100;
    p36_value__105 <= p35_value__105;
    p36_value__106 <= p35_value__106;
    p36_value__109 <= p35_value__109;
    p36_value__112 <= p35_value__112;
    p36_value__115 <= p35_value__115;
    p36_value__118 <= p35_value__118;
  end

  // ===== Pipe stage 37:
  wire [1:0] p37_bit_slice_61588_comb;
  wire [1:0] p37_S0__227_comb;
  wire [10:0] p37_S0__226_comb;
  wire [8:0] p37_S0__225_comb;
  wire [9:0] p37_S0__224_comb;
  wire [31:0] p37_and_61586_comb;
  wire [9:0] p37_s_1__175_comb;
  wire [6:0] p37_s_1__174_comb;
  wire [1:0] p37_s_1__173_comb;
  wire [12:0] p37_s_1__172_comb;
  wire [31:0] p37_S0__41_comb;
  wire [31:0] p37_maj__41_comb;
  wire [31:0] p37_s_1__32_comb;
  wire [31:0] p37_e__42_comb;
  wire [31:0] p37_temp2__41_comb;
  wire [31:0] p37_value__95_comb;
  wire [31:0] p37_a__42_comb;
  wire [31:0] p37_value__96_comb;
  wire [5:0] p37_S1__231_comb;
  wire [4:0] p37_S1__230_comb;
  wire [13:0] p37_S1__229_comb;
  wire [6:0] p37_S1__228_comb;
  wire [27:0] p37_add_61561_comb;
  wire [31:0] p37_S1__42_comb;
  wire [31:0] p37_ch__42_comb;
  wire [31:0] p37_temp1__300_comb;
  wire [1:0] p37_S0__231_comb;
  wire [10:0] p37_S0__230_comb;
  wire [8:0] p37_S0__229_comb;
  wire [9:0] p37_S0__228_comb;
  wire [31:0] p37_and_61609_comb;
  wire [9:0] p37_s_1__183_comb;
  wire [6:0] p37_s_1__182_comb;
  wire [1:0] p37_s_1__181_comb;
  wire [12:0] p37_s_1__180_comb;
  wire [31:0] p37_temp1__383_comb;
  wire [31:0] p37_temp1__384_comb;
  wire [31:0] p37_S0__42_comb;
  wire [31:0] p37_maj__42_comb;
  wire [31:0] p37_s_1__34_comb;
  wire [2:0] p37_s_0__211_comb;
  wire [3:0] p37_s_0__210_comb;
  wire [10:0] p37_s_0__209_comb;
  wire [13:0] p37_s_0__208_comb;
  wire [2:0] p37_s_0__215_comb;
  wire [3:0] p37_s_0__214_comb;
  wire [10:0] p37_s_0__213_comb;
  wire [13:0] p37_s_0__212_comb;
  wire [2:0] p37_s_0__219_comb;
  wire [3:0] p37_s_0__218_comb;
  wire [10:0] p37_s_0__217_comb;
  wire [13:0] p37_s_0__216_comb;
  wire [31:0] p37_temp1__385_comb;
  wire [31:0] p37_temp2__42_comb;
  wire [31:0] p37_value__101_comb;
  wire [31:0] p37_s_0__41_comb;
  wire [31:0] p37_s_0__42_comb;
  wire [31:0] p37_s_0__43_comb;
  wire [31:0] p37_e__43_comb;
  wire [31:0] p37_a__43_comb;
  wire [31:0] p37_value__102_comb;
  wire [31:0] p37_value__121_comb;
  wire [31:0] p37_value__124_comb;
  wire [31:0] p37_value__127_comb;
  assign p37_bit_slice_61588_comb = p36_value__90[1:0];
  assign p37_S0__227_comb = p36_a__41[1:0] ^ p36_a__41[12:11] ^ p36_a__41[21:20];
  assign p37_S0__226_comb = p36_a__41[31:21] ^ p36_a__41[10:0] ^ p36_a__41[19:9];
  assign p37_S0__225_comb = p36_a__41[20:12] ^ p36_a__41[31:23] ^ p36_a__41[8:0];
  assign p37_S0__224_comb = p36_a__41[11:2] ^ p36_a__41[22:13] ^ p36_a__41[31:22];
  assign p37_and_61586_comb = p36_a__41 & p36_a__40;
  assign p37_s_1__175_comb = p36_value__90[16:7] ^ p36_value__90[18:9];
  assign p37_s_1__174_comb = p36_value__90[6:0] ^ p36_value__90[8:2] ^ p36_value__90[31:25];
  assign p37_s_1__173_comb = p36_value__90[31:30] ^ p37_bit_slice_61588_comb ^ p36_value__90[24:23];
  assign p37_s_1__172_comb = p36_value__90[29:17] ^ p36_value__90[31:19] ^ p36_value__90[22:10];
  assign p37_S0__41_comb = {p37_S0__227_comb, p37_S0__226_comb, p37_S0__225_comb, p37_S0__224_comb};
  assign p37_maj__41_comb = p37_and_61586_comb ^ p36_a__41 & p36_a__39 ^ p36_and_61483;
  assign p37_s_1__32_comb = {p37_s_1__175_comb, p37_s_1__174_comb, p37_s_1__173_comb, p37_s_1__172_comb};
  assign p37_e__42_comb = p36_a__38 + p36_temp1__168;
  assign p37_temp2__41_comb = p37_S0__41_comb + p37_maj__41_comb;
  assign p37_value__95_comb = p36_value__75 + p37_s_1__32_comb;
  assign p37_a__42_comb = p36_temp1__168 + p37_temp2__41_comb;
  assign p37_value__96_comb = p36_value__94 + p37_value__95_comb;
  assign p37_S1__231_comb = p37_e__42_comb[5:0] ^ p37_e__42_comb[10:5] ^ p37_e__42_comb[24:19];
  assign p37_S1__230_comb = p37_e__42_comb[31:27] ^ p37_e__42_comb[4:0] ^ p37_e__42_comb[18:14];
  assign p37_S1__229_comb = p37_e__42_comb[26:13] ^ p37_e__42_comb[31:18] ^ p37_e__42_comb[13:0];
  assign p37_S1__228_comb = p37_e__42_comb[12:6] ^ p37_e__42_comb[17:11] ^ p37_e__42_comb[31:25];
  assign p37_add_61561_comb = p36_value__81[31:4] + 28'hc24_b8b7;
  assign p37_S1__42_comb = {p37_S1__231_comb, p37_S1__230_comb, p37_S1__229_comb, p37_S1__228_comb};
  assign p37_ch__42_comb = p37_e__42_comb & p36_e__41 ^ ~(p37_e__42_comb | ~p36_e__40);
  assign p37_temp1__300_comb = {p37_add_61561_comb, p36_value__81[3:0]};
  assign p37_S0__231_comb = p37_a__42_comb[1:0] ^ p37_a__42_comb[12:11] ^ p37_a__42_comb[21:20];
  assign p37_S0__230_comb = p37_a__42_comb[31:21] ^ p37_a__42_comb[10:0] ^ p37_a__42_comb[19:9];
  assign p37_S0__229_comb = p37_a__42_comb[20:12] ^ p37_a__42_comb[31:23] ^ p37_a__42_comb[8:0];
  assign p37_S0__228_comb = p37_a__42_comb[11:2] ^ p37_a__42_comb[22:13] ^ p37_a__42_comb[31:22];
  assign p37_and_61609_comb = p37_a__42_comb & p36_a__41;
  assign p37_s_1__183_comb = p37_value__96_comb[16:7] ^ p37_value__96_comb[18:9];
  assign p37_s_1__182_comb = p37_value__96_comb[6:0] ^ p37_value__96_comb[8:2] ^ p37_value__96_comb[31:25];
  assign p37_s_1__181_comb = p37_value__96_comb[31:30] ^ p37_value__96_comb[1:0] ^ p37_value__96_comb[24:23];
  assign p37_s_1__180_comb = p37_value__96_comb[29:17] ^ p37_value__96_comb[31:19] ^ p37_value__96_comb[22:10];
  assign p37_temp1__383_comb = p36_e__39 + p37_S1__42_comb;
  assign p37_temp1__384_comb = p37_ch__42_comb + p37_temp1__300_comb;
  assign p37_S0__42_comb = {p37_S0__231_comb, p37_S0__230_comb, p37_S0__229_comb, p37_S0__228_comb};
  assign p37_maj__42_comb = p37_and_61609_comb ^ p37_a__42_comb & p36_a__40 ^ p37_and_61586_comb;
  assign p37_s_1__34_comb = {p37_s_1__183_comb, p37_s_1__182_comb, p37_s_1__181_comb, p37_s_1__180_comb};
  assign p37_s_0__211_comb = p36_value__78[6:4] ^ p36_value__78[17:15];
  assign p37_s_0__210_comb = p36_value__78[3:0] ^ p36_value__78[14:11] ^ p36_value__78[31:28];
  assign p37_s_0__209_comb = p36_value__78[31:21] ^ p36_value__78[10:0] ^ p36_value__78[27:17];
  assign p37_s_0__208_comb = p36_value__78[20:7] ^ p36_value__78[31:18] ^ p36_value__78[16:3];
  assign p37_s_0__215_comb = p36_value__81[6:4] ^ p36_value__81[17:15];
  assign p37_s_0__214_comb = p36_value__81[3:0] ^ p36_value__81[14:11] ^ p36_value__81[31:28];
  assign p37_s_0__213_comb = p36_value__81[31:21] ^ p36_value__81[10:0] ^ p36_value__81[27:17];
  assign p37_s_0__212_comb = p36_value__81[20:7] ^ p36_value__81[31:18] ^ p36_value__81[16:3];
  assign p37_s_0__219_comb = p36_value__84[6:4] ^ p36_value__84[17:15];
  assign p37_s_0__218_comb = p36_value__84[3:0] ^ p36_value__84[14:11] ^ p36_value__84[31:28];
  assign p37_s_0__217_comb = p36_value__84[31:21] ^ p36_value__84[10:0] ^ p36_value__84[27:17];
  assign p37_s_0__216_comb = p36_value__84[20:7] ^ p36_value__84[31:18] ^ p36_value__84[16:3];
  assign p37_temp1__385_comb = p37_temp1__383_comb + p37_temp1__384_comb;
  assign p37_temp2__42_comb = p37_S0__42_comb + p37_maj__42_comb;
  assign p37_value__101_comb = p36_value__81 + p37_s_1__34_comb;
  assign p37_s_0__41_comb = {p37_s_0__211_comb, p37_s_0__210_comb, p37_s_0__209_comb, p37_s_0__208_comb};
  assign p37_s_0__42_comb = {p37_s_0__215_comb, p37_s_0__214_comb, p37_s_0__213_comb, p37_s_0__212_comb};
  assign p37_s_0__43_comb = {p37_s_0__219_comb, p37_s_0__218_comb, p37_s_0__217_comb, p37_s_0__216_comb};
  assign p37_e__43_comb = p36_a__39 + p37_temp1__385_comb;
  assign p37_a__43_comb = p37_temp1__385_comb + p37_temp2__42_comb;
  assign p37_value__102_comb = p36_value__100 + p37_value__101_comb;
  assign p37_value__121_comb = p36_value__75 + p37_s_0__41_comb;
  assign p37_value__124_comb = p36_value__78 + p37_s_0__42_comb;
  assign p37_value__127_comb = p36_value__81 + p37_s_0__43_comb;

  // Registers for pipe stage 37:
  reg [31:0] p37_e__40;
  reg [31:0] p37_e__41;
  reg [31:0] p37_e__42;
  reg [31:0] p37_e__43;
  reg [31:0] p37_value__84;
  reg [31:0] p37_a__40;
  reg [31:0] p37_value__87;
  reg [31:0] p37_a__41;
  reg [31:0] p37_value__90;
  reg [1:0] p37_bit_slice_61588;
  reg [31:0] p37_a__42;
  reg [31:0] p37_and_61609;
  reg [31:0] p37_value__93;
  reg [31:0] p37_a__43;
  reg [31:0] p37_value__96;
  reg [31:0] p37_value__99;
  reg [31:0] p37_value__102;
  reg [31:0] p37_value__105;
  reg [31:0] p37_value__106;
  reg [31:0] p37_value__109;
  reg [31:0] p37_value__112;
  reg [31:0] p37_value__115;
  reg [31:0] p37_value__118;
  reg [31:0] p37_value__121;
  reg [31:0] p37_value__124;
  reg [31:0] p37_value__127;
  always_ff @ (posedge clk) begin
    p37_e__40 <= p36_e__40;
    p37_e__41 <= p36_e__41;
    p37_e__42 <= p37_e__42_comb;
    p37_e__43 <= p37_e__43_comb;
    p37_value__84 <= p36_value__84;
    p37_a__40 <= p36_a__40;
    p37_value__87 <= p36_value__87;
    p37_a__41 <= p36_a__41;
    p37_value__90 <= p36_value__90;
    p37_bit_slice_61588 <= p37_bit_slice_61588_comb;
    p37_a__42 <= p37_a__42_comb;
    p37_and_61609 <= p37_and_61609_comb;
    p37_value__93 <= p36_value__93;
    p37_a__43 <= p37_a__43_comb;
    p37_value__96 <= p37_value__96_comb;
    p37_value__99 <= p36_value__99;
    p37_value__102 <= p37_value__102_comb;
    p37_value__105 <= p36_value__105;
    p37_value__106 <= p36_value__106;
    p37_value__109 <= p36_value__109;
    p37_value__112 <= p36_value__112;
    p37_value__115 <= p36_value__115;
    p37_value__118 <= p36_value__118;
    p37_value__121 <= p37_value__121_comb;
    p37_value__124 <= p37_value__124_comb;
    p37_value__127 <= p37_value__127_comb;
  end

  // ===== Pipe stage 38:
  wire [9:0] p38_s_1__191_comb;
  wire [6:0] p38_s_1__190_comb;
  wire [1:0] p38_s_1__189_comb;
  wire [12:0] p38_s_1__188_comb;
  wire [31:0] p38_s_1__36_comb;
  wire [31:0] p38_value__107_comb;
  wire [5:0] p38_S1__235_comb;
  wire [4:0] p38_S1__234_comb;
  wire [13:0] p38_S1__233_comb;
  wire [6:0] p38_S1__232_comb;
  wire [31:0] p38_value__108_comb;
  wire [31:0] p38_S1__43_comb;
  wire [31:0] p38_temp1__173_comb;
  wire [31:0] p38_ch__43_comb;
  wire [1:0] p38_S0__235_comb;
  wire [10:0] p38_S0__234_comb;
  wire [8:0] p38_S0__233_comb;
  wire [9:0] p38_S0__232_comb;
  wire [31:0] p38_and_61795_comb;
  wire [9:0] p38_s_1__199_comb;
  wire [6:0] p38_s_1__198_comb;
  wire [1:0] p38_s_1__197_comb;
  wire [12:0] p38_s_1__196_comb;
  wire [31:0] p38_temp1__174_comb;
  wire [31:0] p38_temp1__301_comb;
  wire [31:0] p38_S0__43_comb;
  wire [31:0] p38_maj__43_comb;
  wire [31:0] p38_s_1__38_comb;
  wire [2:0] p38_s_0__223_comb;
  wire [3:0] p38_s_0__222_comb;
  wire [10:0] p38_s_0__221_comb;
  wire [13:0] p38_s_0__220_comb;
  wire [31:0] p38_temp1__176_comb;
  wire [31:0] p38_temp2__43_comb;
  wire [31:0] p38_value__113_comb;
  wire [31:0] p38_s_0__44_comb;
  wire [31:0] p38_e__44_comb;
  wire [31:0] p38_a__44_comb;
  wire [31:0] p38_value__114_comb;
  wire [31:0] p38_value__130_comb;
  assign p38_s_1__191_comb = p37_value__102[16:7] ^ p37_value__102[18:9];
  assign p38_s_1__190_comb = p37_value__102[6:0] ^ p37_value__102[8:2] ^ p37_value__102[31:25];
  assign p38_s_1__189_comb = p37_value__102[31:30] ^ p37_value__102[1:0] ^ p37_value__102[24:23];
  assign p38_s_1__188_comb = p37_value__102[29:17] ^ p37_value__102[31:19] ^ p37_value__102[22:10];
  assign p38_s_1__36_comb = {p38_s_1__191_comb, p38_s_1__190_comb, p38_s_1__189_comb, p38_s_1__188_comb};
  assign p38_value__107_comb = p37_value__87 + p38_s_1__36_comb;
  assign p38_S1__235_comb = p37_e__43[5:0] ^ p37_e__43[10:5] ^ p37_e__43[24:19];
  assign p38_S1__234_comb = p37_e__43[31:27] ^ p37_e__43[4:0] ^ p37_e__43[18:14];
  assign p38_S1__233_comb = p37_e__43[26:13] ^ p37_e__43[31:18] ^ p37_e__43[13:0];
  assign p38_S1__232_comb = p37_e__43[12:6] ^ p37_e__43[17:11] ^ p37_e__43[31:25];
  assign p38_value__108_comb = p37_value__106 + p38_value__107_comb;
  assign p38_S1__43_comb = {p38_S1__235_comb, p38_S1__234_comb, p38_S1__233_comb, p38_S1__232_comb};
  assign p38_temp1__173_comb = p37_e__40 + p38_S1__43_comb;
  assign p38_ch__43_comb = p37_e__43 & p37_e__42 ^ ~(p37_e__43 | ~p37_e__41);
  assign p38_S0__235_comb = p37_a__43[1:0] ^ p37_a__43[12:11] ^ p37_a__43[21:20];
  assign p38_S0__234_comb = p37_a__43[31:21] ^ p37_a__43[10:0] ^ p37_a__43[19:9];
  assign p38_S0__233_comb = p37_a__43[20:12] ^ p37_a__43[31:23] ^ p37_a__43[8:0];
  assign p38_S0__232_comb = p37_a__43[11:2] ^ p37_a__43[22:13] ^ p37_a__43[31:22];
  assign p38_and_61795_comb = p37_a__43 & p37_a__42;
  assign p38_s_1__199_comb = p38_value__108_comb[16:7] ^ p38_value__108_comb[18:9];
  assign p38_s_1__198_comb = p38_value__108_comb[6:0] ^ p38_value__108_comb[8:2] ^ p38_value__108_comb[31:25];
  assign p38_s_1__197_comb = p38_value__108_comb[31:30] ^ p38_value__108_comb[1:0] ^ p38_value__108_comb[24:23];
  assign p38_s_1__196_comb = p38_value__108_comb[29:17] ^ p38_value__108_comb[31:19] ^ p38_value__108_comb[22:10];
  assign p38_temp1__174_comb = p38_temp1__173_comb + p38_ch__43_comb;
  assign p38_temp1__301_comb = p37_value__84 + 32'hc76c_51a3;
  assign p38_S0__43_comb = {p38_S0__235_comb, p38_S0__234_comb, p38_S0__233_comb, p38_S0__232_comb};
  assign p38_maj__43_comb = p38_and_61795_comb ^ p37_a__43 & p37_a__41 ^ p37_and_61609;
  assign p38_s_1__38_comb = {p38_s_1__199_comb, p38_s_1__198_comb, p38_s_1__197_comb, p38_s_1__196_comb};
  assign p38_s_0__223_comb = p37_value__87[6:4] ^ p37_value__87[17:15];
  assign p38_s_0__222_comb = p37_value__87[3:0] ^ p37_value__87[14:11] ^ p37_value__87[31:28];
  assign p38_s_0__221_comb = p37_value__87[31:21] ^ p37_value__87[10:0] ^ p37_value__87[27:17];
  assign p38_s_0__220_comb = p37_value__87[20:7] ^ p37_value__87[31:18] ^ p37_value__87[16:3];
  assign p38_temp1__176_comb = p38_temp1__174_comb + p38_temp1__301_comb;
  assign p38_temp2__43_comb = p38_S0__43_comb + p38_maj__43_comb;
  assign p38_value__113_comb = p37_value__93 + p38_s_1__38_comb;
  assign p38_s_0__44_comb = {p38_s_0__223_comb, p38_s_0__222_comb, p38_s_0__221_comb, p38_s_0__220_comb};
  assign p38_e__44_comb = p37_a__40 + p38_temp1__176_comb;
  assign p38_a__44_comb = p38_temp1__176_comb + p38_temp2__43_comb;
  assign p38_value__114_comb = p37_value__112 + p38_value__113_comb;
  assign p38_value__130_comb = p37_value__84 + p38_s_0__44_comb;

  // Registers for pipe stage 38:
  reg [31:0] p38_e__41;
  reg [31:0] p38_e__42;
  reg [31:0] p38_e__43;
  reg [31:0] p38_e__44;
  reg [31:0] p38_value__87;
  reg [31:0] p38_a__41;
  reg [31:0] p38_value__90;
  reg [1:0] p38_bit_slice_61588;
  reg [31:0] p38_a__42;
  reg [31:0] p38_value__93;
  reg [31:0] p38_a__43;
  reg [31:0] p38_value__96;
  reg [31:0] p38_and_61795;
  reg [31:0] p38_a__44;
  reg [31:0] p38_value__99;
  reg [31:0] p38_value__102;
  reg [31:0] p38_value__105;
  reg [31:0] p38_value__108;
  reg [31:0] p38_value__109;
  reg [31:0] p38_value__114;
  reg [31:0] p38_value__115;
  reg [31:0] p38_value__118;
  reg [31:0] p38_value__121;
  reg [31:0] p38_value__124;
  reg [31:0] p38_value__127;
  reg [31:0] p38_value__130;
  always_ff @ (posedge clk) begin
    p38_e__41 <= p37_e__41;
    p38_e__42 <= p37_e__42;
    p38_e__43 <= p37_e__43;
    p38_e__44 <= p38_e__44_comb;
    p38_value__87 <= p37_value__87;
    p38_a__41 <= p37_a__41;
    p38_value__90 <= p37_value__90;
    p38_bit_slice_61588 <= p37_bit_slice_61588;
    p38_a__42 <= p37_a__42;
    p38_value__93 <= p37_value__93;
    p38_a__43 <= p37_a__43;
    p38_value__96 <= p37_value__96;
    p38_and_61795 <= p38_and_61795_comb;
    p38_a__44 <= p38_a__44_comb;
    p38_value__99 <= p37_value__99;
    p38_value__102 <= p37_value__102;
    p38_value__105 <= p37_value__105;
    p38_value__108 <= p38_value__108_comb;
    p38_value__109 <= p37_value__109;
    p38_value__114 <= p38_value__114_comb;
    p38_value__115 <= p37_value__115;
    p38_value__118 <= p37_value__118;
    p38_value__121 <= p37_value__121;
    p38_value__124 <= p37_value__124;
    p38_value__127 <= p37_value__127;
    p38_value__130 <= p38_value__130_comb;
  end

  // ===== Pipe stage 39:
  wire [9:0] p39_s_1__195_comb;
  wire [6:0] p39_s_1__194_comb;
  wire [1:0] p39_s_1__193_comb;
  wire [12:0] p39_s_1__192_comb;
  wire [9:0] p39_s_1__207_comb;
  wire [6:0] p39_s_1__206_comb;
  wire [1:0] p39_s_1__205_comb;
  wire [12:0] p39_s_1__204_comb;
  wire [31:0] p39_s_1__37_comb;
  wire [31:0] p39_s_1__40_comb;
  wire [31:0] p39_value__110_comb;
  wire [31:0] p39_value__119_comb;
  wire [5:0] p39_S1__239_comb;
  wire [4:0] p39_S1__238_comb;
  wire [13:0] p39_S1__237_comb;
  wire [6:0] p39_S1__236_comb;
  wire [31:0] p39_value__111_comb;
  wire [31:0] p39_value__120_comb;
  wire [31:0] p39_S1__44_comb;
  wire [31:0] p39_temp1__177_comb;
  wire [31:0] p39_ch__44_comb;
  wire [1:0] p39_S0__239_comb;
  wire [10:0] p39_S0__238_comb;
  wire [8:0] p39_S0__237_comb;
  wire [9:0] p39_S0__236_comb;
  wire [31:0] p39_and_61953_comb;
  wire [9:0] p39_s_1__203_comb;
  wire [6:0] p39_s_1__202_comb;
  wire [1:0] p39_s_1__201_comb;
  wire [12:0] p39_s_1__200_comb;
  wire [9:0] p39_s_1__215_comb;
  wire [6:0] p39_s_1__214_comb;
  wire [1:0] p39_s_1__213_comb;
  wire [12:0] p39_s_1__212_comb;
  wire [31:0] p39_temp1__178_comb;
  wire [31:0] p39_temp1__302_comb;
  wire [31:0] p39_S0__44_comb;
  wire [31:0] p39_maj__44_comb;
  wire [31:0] p39_s_1__39_comb;
  wire [31:0] p39_s_1__42_comb;
  wire [2:0] p39_s_0__227_comb;
  wire [3:0] p39_s_0__226_comb;
  wire [10:0] p39_s_0__225_comb;
  wire [13:0] p39_s_0__224_comb;
  wire [2:0] p39_s_0__231_comb;
  wire [3:0] p39_s_0__230_comb;
  wire [10:0] p39_s_0__229_comb;
  wire [13:0] p39_s_0__228_comb;
  wire [31:0] p39_temp1__180_comb;
  wire [29:0] p39_add_61935_comb;
  wire [31:0] p39_temp2__44_comb;
  wire [29:0] p39_add_61961_comb;
  wire [31:0] p39_value__116_comb;
  wire [31:0] p39_value__125_comb;
  wire [31:0] p39_s_0__45_comb;
  wire [31:0] p39_s_0__46_comb;
  wire [31:0] p39_e__45_comb;
  wire [31:0] p39_temp1__303_comb;
  wire [31:0] p39_a__45_comb;
  wire [31:0] p39_temp1__308_comb;
  wire [31:0] p39_value__117_comb;
  wire [31:0] p39_value__126_comb;
  wire [31:0] p39_value__133_comb;
  wire [31:0] p39_value__136_comb;
  assign p39_s_1__195_comb = p38_value__105[16:7] ^ p38_value__105[18:9];
  assign p39_s_1__194_comb = p38_value__105[6:0] ^ p38_value__105[8:2] ^ p38_value__105[31:25];
  assign p39_s_1__193_comb = p38_value__105[31:30] ^ p38_value__105[1:0] ^ p38_value__105[24:23];
  assign p39_s_1__192_comb = p38_value__105[29:17] ^ p38_value__105[31:19] ^ p38_value__105[22:10];
  assign p39_s_1__207_comb = p38_value__114[16:7] ^ p38_value__114[18:9];
  assign p39_s_1__206_comb = p38_value__114[6:0] ^ p38_value__114[8:2] ^ p38_value__114[31:25];
  assign p39_s_1__205_comb = p38_value__114[31:30] ^ p38_value__114[1:0] ^ p38_value__114[24:23];
  assign p39_s_1__204_comb = p38_value__114[29:17] ^ p38_value__114[31:19] ^ p38_value__114[22:10];
  assign p39_s_1__37_comb = {p39_s_1__195_comb, p39_s_1__194_comb, p39_s_1__193_comb, p39_s_1__192_comb};
  assign p39_s_1__40_comb = {p39_s_1__207_comb, p39_s_1__206_comb, p39_s_1__205_comb, p39_s_1__204_comb};
  assign p39_value__110_comb = p38_value__90 + p39_s_1__37_comb;
  assign p39_value__119_comb = p38_value__99 + p39_s_1__40_comb;
  assign p39_S1__239_comb = p38_e__44[5:0] ^ p38_e__44[10:5] ^ p38_e__44[24:19];
  assign p39_S1__238_comb = p38_e__44[31:27] ^ p38_e__44[4:0] ^ p38_e__44[18:14];
  assign p39_S1__237_comb = p38_e__44[26:13] ^ p38_e__44[31:18] ^ p38_e__44[13:0];
  assign p39_S1__236_comb = p38_e__44[12:6] ^ p38_e__44[17:11] ^ p38_e__44[31:25];
  assign p39_value__111_comb = p38_value__109 + p39_value__110_comb;
  assign p39_value__120_comb = p38_value__118 + p39_value__119_comb;
  assign p39_S1__44_comb = {p39_S1__239_comb, p39_S1__238_comb, p39_S1__237_comb, p39_S1__236_comb};
  assign p39_temp1__177_comb = p38_e__41 + p39_S1__44_comb;
  assign p39_ch__44_comb = p38_e__44 & p38_e__43 ^ ~(p38_e__44 | ~p38_e__42);
  assign p39_S0__239_comb = p38_a__44[1:0] ^ p38_a__44[12:11] ^ p38_a__44[21:20];
  assign p39_S0__238_comb = p38_a__44[31:21] ^ p38_a__44[10:0] ^ p38_a__44[19:9];
  assign p39_S0__237_comb = p38_a__44[20:12] ^ p38_a__44[31:23] ^ p38_a__44[8:0];
  assign p39_S0__236_comb = p38_a__44[11:2] ^ p38_a__44[22:13] ^ p38_a__44[31:22];
  assign p39_and_61953_comb = p38_a__44 & p38_a__43;
  assign p39_s_1__203_comb = p39_value__111_comb[16:7] ^ p39_value__111_comb[18:9];
  assign p39_s_1__202_comb = p39_value__111_comb[6:0] ^ p39_value__111_comb[8:2] ^ p39_value__111_comb[31:25];
  assign p39_s_1__201_comb = p39_value__111_comb[31:30] ^ p39_value__111_comb[1:0] ^ p39_value__111_comb[24:23];
  assign p39_s_1__200_comb = p39_value__111_comb[29:17] ^ p39_value__111_comb[31:19] ^ p39_value__111_comb[22:10];
  assign p39_s_1__215_comb = p39_value__120_comb[16:7] ^ p39_value__120_comb[18:9];
  assign p39_s_1__214_comb = p39_value__120_comb[6:0] ^ p39_value__120_comb[8:2] ^ p39_value__120_comb[31:25];
  assign p39_s_1__213_comb = p39_value__120_comb[31:30] ^ p39_value__120_comb[1:0] ^ p39_value__120_comb[24:23];
  assign p39_s_1__212_comb = p39_value__120_comb[29:17] ^ p39_value__120_comb[31:19] ^ p39_value__120_comb[22:10];
  assign p39_temp1__178_comb = p39_temp1__177_comb + p39_ch__44_comb;
  assign p39_temp1__302_comb = p38_value__87 + 32'hd192_e819;
  assign p39_S0__44_comb = {p39_S0__239_comb, p39_S0__238_comb, p39_S0__237_comb, p39_S0__236_comb};
  assign p39_maj__44_comb = p39_and_61953_comb ^ p38_a__44 & p38_a__42 ^ p38_and_61795;
  assign p39_s_1__39_comb = {p39_s_1__203_comb, p39_s_1__202_comb, p39_s_1__201_comb, p39_s_1__200_comb};
  assign p39_s_1__42_comb = {p39_s_1__215_comb, p39_s_1__214_comb, p39_s_1__213_comb, p39_s_1__212_comb};
  assign p39_s_0__227_comb = p38_value__90[6:4] ^ p38_value__90[17:15];
  assign p39_s_0__226_comb = p38_value__90[3:0] ^ p38_value__90[14:11] ^ p38_value__90[31:28];
  assign p39_s_0__225_comb = p38_value__90[31:21] ^ p38_value__90[10:0] ^ p38_value__90[27:17];
  assign p39_s_0__224_comb = p38_value__90[20:7] ^ p38_value__90[31:18] ^ p38_value__90[16:3];
  assign p39_s_0__231_comb = p38_value__93[6:4] ^ p38_value__93[17:15];
  assign p39_s_0__230_comb = p38_value__93[3:0] ^ p38_value__93[14:11] ^ p38_value__93[31:28];
  assign p39_s_0__229_comb = p38_value__93[31:21] ^ p38_value__93[10:0] ^ p38_value__93[27:17];
  assign p39_s_0__228_comb = p38_value__93[20:7] ^ p38_value__93[31:18] ^ p38_value__93[16:3];
  assign p39_temp1__180_comb = p39_temp1__178_comb + p39_temp1__302_comb;
  assign p39_add_61935_comb = p38_value__90[31:2] + 30'h35a6_4189;
  assign p39_temp2__44_comb = p39_S0__44_comb + p39_maj__44_comb;
  assign p39_add_61961_comb = p38_value__105[31:2] + 30'h09d2_1dd3;
  assign p39_value__116_comb = p38_value__96 + p39_s_1__39_comb;
  assign p39_value__125_comb = p38_value__105 + p39_s_1__42_comb;
  assign p39_s_0__45_comb = {p39_s_0__227_comb, p39_s_0__226_comb, p39_s_0__225_comb, p39_s_0__224_comb};
  assign p39_s_0__46_comb = {p39_s_0__231_comb, p39_s_0__230_comb, p39_s_0__229_comb, p39_s_0__228_comb};
  assign p39_e__45_comb = p38_a__41 + p39_temp1__180_comb;
  assign p39_temp1__303_comb = {p39_add_61935_comb, p38_bit_slice_61588};
  assign p39_a__45_comb = p39_temp1__180_comb + p39_temp2__44_comb;
  assign p39_temp1__308_comb = {p39_add_61961_comb, p38_value__105[1:0]};
  assign p39_value__117_comb = p38_value__115 + p39_value__116_comb;
  assign p39_value__126_comb = p38_value__124 + p39_value__125_comb;
  assign p39_value__133_comb = p38_value__87 + p39_s_0__45_comb;
  assign p39_value__136_comb = p38_value__90 + p39_s_0__46_comb;

  // Registers for pipe stage 39:
  reg [31:0] p39_e__42;
  reg [31:0] p39_e__43;
  reg [31:0] p39_e__44;
  reg [31:0] p39_e__45;
  reg [31:0] p39_temp1__303;
  reg [31:0] p39_a__42;
  reg [31:0] p39_value__93;
  reg [31:0] p39_a__43;
  reg [31:0] p39_value__96;
  reg [31:0] p39_a__44;
  reg [31:0] p39_value__99;
  reg [31:0] p39_and_61953;
  reg [31:0] p39_a__45;
  reg [31:0] p39_value__102;
  reg [31:0] p39_temp1__308;
  reg [31:0] p39_value__108;
  reg [31:0] p39_value__111;
  reg [31:0] p39_value__114;
  reg [31:0] p39_value__117;
  reg [31:0] p39_value__120;
  reg [31:0] p39_value__121;
  reg [31:0] p39_value__126;
  reg [31:0] p39_value__127;
  reg [31:0] p39_value__130;
  reg [31:0] p39_value__133;
  reg [31:0] p39_value__136;
  always_ff @ (posedge clk) begin
    p39_e__42 <= p38_e__42;
    p39_e__43 <= p38_e__43;
    p39_e__44 <= p38_e__44;
    p39_e__45 <= p39_e__45_comb;
    p39_temp1__303 <= p39_temp1__303_comb;
    p39_a__42 <= p38_a__42;
    p39_value__93 <= p38_value__93;
    p39_a__43 <= p38_a__43;
    p39_value__96 <= p38_value__96;
    p39_a__44 <= p38_a__44;
    p39_value__99 <= p38_value__99;
    p39_and_61953 <= p39_and_61953_comb;
    p39_a__45 <= p39_a__45_comb;
    p39_value__102 <= p38_value__102;
    p39_temp1__308 <= p39_temp1__308_comb;
    p39_value__108 <= p38_value__108;
    p39_value__111 <= p39_value__111_comb;
    p39_value__114 <= p38_value__114;
    p39_value__117 <= p39_value__117_comb;
    p39_value__120 <= p39_value__120_comb;
    p39_value__121 <= p38_value__121;
    p39_value__126 <= p39_value__126_comb;
    p39_value__127 <= p38_value__127;
    p39_value__130 <= p38_value__130;
    p39_value__133 <= p39_value__133_comb;
    p39_value__136 <= p39_value__136_comb;
  end

  // ===== Pipe stage 40:
  wire [5:0] p40_S1__243_comb;
  wire [4:0] p40_S1__242_comb;
  wire [13:0] p40_S1__241_comb;
  wire [6:0] p40_S1__240_comb;
  wire [9:0] p40_s_1__211_comb;
  wire [6:0] p40_s_1__210_comb;
  wire [1:0] p40_s_1__209_comb;
  wire [12:0] p40_s_1__208_comb;
  wire [9:0] p40_s_1__223_comb;
  wire [6:0] p40_s_1__222_comb;
  wire [1:0] p40_s_1__221_comb;
  wire [12:0] p40_s_1__220_comb;
  wire [31:0] p40_S1__45_comb;
  wire [31:0] p40_ch__45_comb;
  wire [31:0] p40_s_1__41_comb;
  wire [31:0] p40_s_1__44_comb;
  wire [31:0] p40_temp1__380_comb;
  wire [31:0] p40_temp1__381_comb;
  wire [31:0] p40_value__122_comb;
  wire [31:0] p40_value__131_comb;
  wire [31:0] p40_temp1__382_comb;
  wire [31:0] p40_value__123_comb;
  wire [31:0] p40_value__132_comb;
  wire [31:0] p40_e__46_comb;
  wire [1:0] p40_S0__243_comb;
  wire [10:0] p40_S0__242_comb;
  wire [8:0] p40_S0__241_comb;
  wire [9:0] p40_S0__240_comb;
  wire [31:0] p40_and_62182_comb;
  wire [9:0] p40_s_1__219_comb;
  wire [6:0] p40_s_1__218_comb;
  wire [1:0] p40_s_1__217_comb;
  wire [12:0] p40_s_1__216_comb;
  wire [9:0] p40_s_1__231_comb;
  wire [6:0] p40_s_1__230_comb;
  wire [1:0] p40_s_1__229_comb;
  wire [12:0] p40_s_1__228_comb;
  wire [5:0] p40_S1__247_comb;
  wire [4:0] p40_S1__246_comb;
  wire [13:0] p40_S1__245_comb;
  wire [6:0] p40_S1__244_comb;
  wire [31:0] p40_S0__45_comb;
  wire [31:0] p40_maj__45_comb;
  wire [31:0] p40_s_1__43_comb;
  wire [31:0] p40_s_1__46_comb;
  wire [31:0] p40_S1__46_comb;
  wire [28:0] p40_add_62184_comb;
  wire [31:0] p40_temp2__45_comb;
  wire [31:0] p40_value__128_comb;
  wire [28:0] p40_add_62255_comb;
  wire [31:0] p40_value__137_comb;
  wire [31:0] p40_temp1__185_comb;
  wire [31:0] p40_temp1__307_comb;
  wire [31:0] p40_a__46_comb;
  wire [31:0] p40_temp1__309_comb;
  wire [31:0] p40_temp1__310_comb;
  wire [31:0] p40_temp1__312_comb;
  wire [31:0] p40_temp1__315_comb;
  wire [31:0] p40_value__129_comb;
  wire [31:0] p40_temp1__317_comb;
  wire [31:0] p40_value__138_comb;
  assign p40_S1__243_comb = p39_e__45[5:0] ^ p39_e__45[10:5] ^ p39_e__45[24:19];
  assign p40_S1__242_comb = p39_e__45[31:27] ^ p39_e__45[4:0] ^ p39_e__45[18:14];
  assign p40_S1__241_comb = p39_e__45[26:13] ^ p39_e__45[31:18] ^ p39_e__45[13:0];
  assign p40_S1__240_comb = p39_e__45[12:6] ^ p39_e__45[17:11] ^ p39_e__45[31:25];
  assign p40_s_1__211_comb = p39_value__117[16:7] ^ p39_value__117[18:9];
  assign p40_s_1__210_comb = p39_value__117[6:0] ^ p39_value__117[8:2] ^ p39_value__117[31:25];
  assign p40_s_1__209_comb = p39_value__117[31:30] ^ p39_value__117[1:0] ^ p39_value__117[24:23];
  assign p40_s_1__208_comb = p39_value__117[29:17] ^ p39_value__117[31:19] ^ p39_value__117[22:10];
  assign p40_s_1__223_comb = p39_value__126[16:7] ^ p39_value__126[18:9];
  assign p40_s_1__222_comb = p39_value__126[6:0] ^ p39_value__126[8:2] ^ p39_value__126[31:25];
  assign p40_s_1__221_comb = p39_value__126[31:30] ^ p39_value__126[1:0] ^ p39_value__126[24:23];
  assign p40_s_1__220_comb = p39_value__126[29:17] ^ p39_value__126[31:19] ^ p39_value__126[22:10];
  assign p40_S1__45_comb = {p40_S1__243_comb, p40_S1__242_comb, p40_S1__241_comb, p40_S1__240_comb};
  assign p40_ch__45_comb = p39_e__45 & p39_e__44 ^ ~(p39_e__45 | ~p39_e__43);
  assign p40_s_1__41_comb = {p40_s_1__211_comb, p40_s_1__210_comb, p40_s_1__209_comb, p40_s_1__208_comb};
  assign p40_s_1__44_comb = {p40_s_1__223_comb, p40_s_1__222_comb, p40_s_1__221_comb, p40_s_1__220_comb};
  assign p40_temp1__380_comb = p39_e__42 + p40_S1__45_comb;
  assign p40_temp1__381_comb = p40_ch__45_comb + p39_temp1__303;
  assign p40_value__122_comb = p39_value__102 + p40_s_1__41_comb;
  assign p40_value__131_comb = p39_value__111 + p40_s_1__44_comb;
  assign p40_temp1__382_comb = p40_temp1__380_comb + p40_temp1__381_comb;
  assign p40_value__123_comb = p39_value__121 + p40_value__122_comb;
  assign p40_value__132_comb = p39_value__130 + p40_value__131_comb;
  assign p40_e__46_comb = p39_a__42 + p40_temp1__382_comb;
  assign p40_S0__243_comb = p39_a__45[1:0] ^ p39_a__45[12:11] ^ p39_a__45[21:20];
  assign p40_S0__242_comb = p39_a__45[31:21] ^ p39_a__45[10:0] ^ p39_a__45[19:9];
  assign p40_S0__241_comb = p39_a__45[20:12] ^ p39_a__45[31:23] ^ p39_a__45[8:0];
  assign p40_S0__240_comb = p39_a__45[11:2] ^ p39_a__45[22:13] ^ p39_a__45[31:22];
  assign p40_and_62182_comb = p39_a__45 & p39_a__44;
  assign p40_s_1__219_comb = p40_value__123_comb[16:7] ^ p40_value__123_comb[18:9];
  assign p40_s_1__218_comb = p40_value__123_comb[6:0] ^ p40_value__123_comb[8:2] ^ p40_value__123_comb[31:25];
  assign p40_s_1__217_comb = p40_value__123_comb[31:30] ^ p40_value__123_comb[1:0] ^ p40_value__123_comb[24:23];
  assign p40_s_1__216_comb = p40_value__123_comb[29:17] ^ p40_value__123_comb[31:19] ^ p40_value__123_comb[22:10];
  assign p40_s_1__231_comb = p40_value__132_comb[16:7] ^ p40_value__132_comb[18:9];
  assign p40_s_1__230_comb = p40_value__132_comb[6:0] ^ p40_value__132_comb[8:2] ^ p40_value__132_comb[31:25];
  assign p40_s_1__229_comb = p40_value__132_comb[31:30] ^ p40_value__132_comb[1:0] ^ p40_value__132_comb[24:23];
  assign p40_s_1__228_comb = p40_value__132_comb[29:17] ^ p40_value__132_comb[31:19] ^ p40_value__132_comb[22:10];
  assign p40_S1__247_comb = p40_e__46_comb[5:0] ^ p40_e__46_comb[10:5] ^ p40_e__46_comb[24:19];
  assign p40_S1__246_comb = p40_e__46_comb[31:27] ^ p40_e__46_comb[4:0] ^ p40_e__46_comb[18:14];
  assign p40_S1__245_comb = p40_e__46_comb[26:13] ^ p40_e__46_comb[31:18] ^ p40_e__46_comb[13:0];
  assign p40_S1__244_comb = p40_e__46_comb[12:6] ^ p40_e__46_comb[17:11] ^ p40_e__46_comb[31:25];
  assign p40_S0__45_comb = {p40_S0__243_comb, p40_S0__242_comb, p40_S0__241_comb, p40_S0__240_comb};
  assign p40_maj__45_comb = p40_and_62182_comb ^ p39_a__45 & p39_a__43 ^ p39_and_61953;
  assign p40_s_1__43_comb = {p40_s_1__219_comb, p40_s_1__218_comb, p40_s_1__217_comb, p40_s_1__216_comb};
  assign p40_s_1__46_comb = {p40_s_1__231_comb, p40_s_1__230_comb, p40_s_1__229_comb, p40_s_1__228_comb};
  assign p40_S1__46_comb = {p40_S1__247_comb, p40_S1__246_comb, p40_S1__245_comb, p40_S1__244_comb};
  assign p40_add_62184_comb = p39_value__102[31:3] + 29'h03c6_ed81;
  assign p40_temp2__45_comb = p40_S0__45_comb + p40_maj__45_comb;
  assign p40_value__128_comb = p39_value__108 + p40_s_1__43_comb;
  assign p40_add_62255_comb = p40_value__132_comb[31:3] + 29'h1198_e041;
  assign p40_value__137_comb = p39_value__117 + p40_s_1__46_comb;
  assign p40_temp1__185_comb = p39_e__43 + p40_S1__46_comb;
  assign p40_temp1__307_comb = {p40_add_62184_comb, p39_value__102[2:0]};
  assign p40_a__46_comb = p40_temp1__382_comb + p40_temp2__45_comb;
  assign p40_temp1__309_comb = p39_value__108 + 32'h34b0_bcb5;
  assign p40_temp1__310_comb = p39_value__111 + 32'h391c_0cb3;
  assign p40_temp1__312_comb = p39_value__117 + 32'h5b9c_ca4f;
  assign p40_temp1__315_comb = p39_value__126 + 32'h78a5_636f;
  assign p40_value__129_comb = p39_value__127 + p40_value__128_comb;
  assign p40_temp1__317_comb = {p40_add_62255_comb, p40_value__132_comb[2:0]};
  assign p40_value__138_comb = p39_value__136 + p40_value__137_comb;

  // Registers for pipe stage 40:
  reg [31:0] p40_e__44;
  reg [31:0] p40_e__45;
  reg [31:0] p40_e__46;
  reg [31:0] p40_temp1__185;
  reg [31:0] p40_value__93;
  reg [31:0] p40_a__43;
  reg [31:0] p40_value__96;
  reg [31:0] p40_a__44;
  reg [31:0] p40_value__99;
  reg [31:0] p40_a__45;
  reg [31:0] p40_and_62182;
  reg [31:0] p40_temp1__307;
  reg [31:0] p40_a__46;
  reg [31:0] p40_temp1__308;
  reg [31:0] p40_temp1__309;
  reg [31:0] p40_temp1__310;
  reg [31:0] p40_value__114;
  reg [31:0] p40_temp1__312;
  reg [31:0] p40_value__120;
  reg [31:0] p40_value__123;
  reg [31:0] p40_temp1__315;
  reg [31:0] p40_value__129;
  reg [31:0] p40_temp1__317;
  reg [31:0] p40_value__133;
  reg [31:0] p40_value__138;
  always_ff @ (posedge clk) begin
    p40_e__44 <= p39_e__44;
    p40_e__45 <= p39_e__45;
    p40_e__46 <= p40_e__46_comb;
    p40_temp1__185 <= p40_temp1__185_comb;
    p40_value__93 <= p39_value__93;
    p40_a__43 <= p39_a__43;
    p40_value__96 <= p39_value__96;
    p40_a__44 <= p39_a__44;
    p40_value__99 <= p39_value__99;
    p40_a__45 <= p39_a__45;
    p40_and_62182 <= p40_and_62182_comb;
    p40_temp1__307 <= p40_temp1__307_comb;
    p40_a__46 <= p40_a__46_comb;
    p40_temp1__308 <= p39_temp1__308;
    p40_temp1__309 <= p40_temp1__309_comb;
    p40_temp1__310 <= p40_temp1__310_comb;
    p40_value__114 <= p39_value__114;
    p40_temp1__312 <= p40_temp1__312_comb;
    p40_value__120 <= p39_value__120;
    p40_value__123 <= p40_value__123_comb;
    p40_temp1__315 <= p40_temp1__315_comb;
    p40_value__129 <= p40_value__129_comb;
    p40_temp1__317 <= p40_temp1__317_comb;
    p40_value__133 <= p39_value__133;
    p40_value__138 <= p40_value__138_comb;
  end

  // ===== Pipe stage 41:
  wire [31:0] p41_ch__46_comb;
  wire [31:0] p41_temp1__186_comb;
  wire [31:0] p41_temp1__304_comb;
  wire [31:0] p41_temp1__188_comb;
  wire [31:0] p41_e__47_comb;
  wire [1:0] p41_S0__247_comb;
  wire [10:0] p41_S0__246_comb;
  wire [8:0] p41_S0__245_comb;
  wire [9:0] p41_S0__244_comb;
  wire [31:0] p41_and_62379_comb;
  wire [9:0] p41_s_1__227_comb;
  wire [6:0] p41_s_1__226_comb;
  wire [1:0] p41_s_1__225_comb;
  wire [12:0] p41_s_1__224_comb;
  wire [5:0] p41_S1__251_comb;
  wire [4:0] p41_S1__250_comb;
  wire [13:0] p41_S1__249_comb;
  wire [6:0] p41_S1__248_comb;
  wire [27:0] p41_add_62356_comb;
  wire [31:0] p41_S0__46_comb;
  wire [31:0] p41_maj__46_comb;
  wire [31:0] p41_s_1__45_comb;
  wire [31:0] p41_S1__47_comb;
  wire [31:0] p41_ch__47_comb;
  wire [31:0] p41_temp1__305_comb;
  wire [31:0] p41_temp2__46_comb;
  wire [30:0] p41_add_62387_comb;
  wire [29:0] p41_add_62392_comb;
  wire [31:0] p41_value__134_comb;
  wire [31:0] p41_temp1__377_comb;
  wire [31:0] p41_temp1__378_comb;
  wire [31:0] p41_a__47_comb;
  wire [31:0] p41_temp1__311_comb;
  wire [31:0] p41_temp1__316_comb;
  wire [31:0] p41_value__135_comb;
  wire [3:0] p41_s_0__234_comb;
  assign p41_ch__46_comb = p40_e__46 & p40_e__45 ^ ~(p40_e__46 | ~p40_e__44);
  assign p41_temp1__186_comb = p40_temp1__185 + p41_ch__46_comb;
  assign p41_temp1__304_comb = p40_value__93 + 32'hf40e_3585;
  assign p41_temp1__188_comb = p41_temp1__186_comb + p41_temp1__304_comb;
  assign p41_e__47_comb = p40_a__43 + p41_temp1__188_comb;
  assign p41_S0__247_comb = p40_a__46[1:0] ^ p40_a__46[12:11] ^ p40_a__46[21:20];
  assign p41_S0__246_comb = p40_a__46[31:21] ^ p40_a__46[10:0] ^ p40_a__46[19:9];
  assign p41_S0__245_comb = p40_a__46[20:12] ^ p40_a__46[31:23] ^ p40_a__46[8:0];
  assign p41_S0__244_comb = p40_a__46[11:2] ^ p40_a__46[22:13] ^ p40_a__46[31:22];
  assign p41_and_62379_comb = p40_a__46 & p40_a__45;
  assign p41_s_1__227_comb = p40_value__129[16:7] ^ p40_value__129[18:9];
  assign p41_s_1__226_comb = p40_value__129[6:0] ^ p40_value__129[8:2] ^ p40_value__129[31:25];
  assign p41_s_1__225_comb = p40_value__129[31:30] ^ p40_value__129[1:0] ^ p40_value__129[24:23];
  assign p41_s_1__224_comb = p40_value__129[29:17] ^ p40_value__129[31:19] ^ p40_value__129[22:10];
  assign p41_S1__251_comb = p41_e__47_comb[5:0] ^ p41_e__47_comb[10:5] ^ p41_e__47_comb[24:19];
  assign p41_S1__250_comb = p41_e__47_comb[31:27] ^ p41_e__47_comb[4:0] ^ p41_e__47_comb[18:14];
  assign p41_S1__249_comb = p41_e__47_comb[26:13] ^ p41_e__47_comb[31:18] ^ p41_e__47_comb[13:0];
  assign p41_S1__248_comb = p41_e__47_comb[12:6] ^ p41_e__47_comb[17:11] ^ p41_e__47_comb[31:25];
  assign p41_add_62356_comb = p40_value__96[31:4] + 28'h106_aa07;
  assign p41_S0__46_comb = {p41_S0__247_comb, p41_S0__246_comb, p41_S0__245_comb, p41_S0__244_comb};
  assign p41_maj__46_comb = p41_and_62379_comb ^ p40_a__46 & p40_a__44 ^ p40_and_62182;
  assign p41_s_1__45_comb = {p41_s_1__227_comb, p41_s_1__226_comb, p41_s_1__225_comb, p41_s_1__224_comb};
  assign p41_S1__47_comb = {p41_S1__251_comb, p41_S1__250_comb, p41_S1__249_comb, p41_S1__248_comb};
  assign p41_ch__47_comb = p41_e__47_comb & p40_e__46 ^ ~(p41_e__47_comb | ~p40_e__45);
  assign p41_temp1__305_comb = {p41_add_62356_comb, p40_value__96[3:0]};
  assign p41_temp2__46_comb = p41_S0__46_comb + p41_maj__46_comb;
  assign p41_add_62387_comb = p40_value__114[31:1] + 31'h276c_5525;
  assign p41_add_62392_comb = p40_value__129[31:2] + 30'h2132_1e05;
  assign p41_value__134_comb = p40_value__114 + p41_s_1__45_comb;
  assign p41_temp1__377_comb = p40_e__44 + p41_S1__47_comb;
  assign p41_temp1__378_comb = p41_ch__47_comb + p41_temp1__305_comb;
  assign p41_a__47_comb = p41_temp1__188_comb + p41_temp2__46_comb;
  assign p41_temp1__311_comb = {p41_add_62387_comb, p40_value__114[0]};
  assign p41_temp1__316_comb = {p41_add_62392_comb, p40_value__129[1:0]};
  assign p41_value__135_comb = p40_value__133 + p41_value__134_comb;
  assign p41_s_0__234_comb = p40_value__96[3:0] ^ p40_value__96[14:11] ^ p40_value__96[31:28];

  // Registers for pipe stage 41:
  reg [31:0] p41_e__45;
  reg [31:0] p41_e__46;
  reg [31:0] p41_value__93;
  reg [31:0] p41_e__47;
  reg [31:0] p41_value__96;
  reg [31:0] p41_temp1__377;
  reg [31:0] p41_temp1__378;
  reg [31:0] p41_a__44;
  reg [31:0] p41_value__99;
  reg [31:0] p41_a__45;
  reg [31:0] p41_temp1__307;
  reg [31:0] p41_a__46;
  reg [31:0] p41_and_62379;
  reg [31:0] p41_temp1__308;
  reg [31:0] p41_a__47;
  reg [31:0] p41_temp1__309;
  reg [31:0] p41_temp1__310;
  reg [31:0] p41_temp1__311;
  reg [31:0] p41_temp1__312;
  reg [31:0] p41_value__120;
  reg [31:0] p41_value__123;
  reg [31:0] p41_temp1__315;
  reg [31:0] p41_temp1__316;
  reg [31:0] p41_temp1__317;
  reg [31:0] p41_value__135;
  reg [31:0] p41_value__138;
  reg [3:0] p41_s_0__234;
  always_ff @ (posedge clk) begin
    p41_e__45 <= p40_e__45;
    p41_e__46 <= p40_e__46;
    p41_value__93 <= p40_value__93;
    p41_e__47 <= p41_e__47_comb;
    p41_value__96 <= p40_value__96;
    p41_temp1__377 <= p41_temp1__377_comb;
    p41_temp1__378 <= p41_temp1__378_comb;
    p41_a__44 <= p40_a__44;
    p41_value__99 <= p40_value__99;
    p41_a__45 <= p40_a__45;
    p41_temp1__307 <= p40_temp1__307;
    p41_a__46 <= p40_a__46;
    p41_and_62379 <= p41_and_62379_comb;
    p41_temp1__308 <= p40_temp1__308;
    p41_a__47 <= p41_a__47_comb;
    p41_temp1__309 <= p40_temp1__309;
    p41_temp1__310 <= p40_temp1__310;
    p41_temp1__311 <= p41_temp1__311_comb;
    p41_temp1__312 <= p40_temp1__312;
    p41_value__120 <= p40_value__120;
    p41_value__123 <= p40_value__123;
    p41_temp1__315 <= p40_temp1__315;
    p41_temp1__316 <= p41_temp1__316_comb;
    p41_temp1__317 <= p40_temp1__317;
    p41_value__135 <= p41_value__135_comb;
    p41_value__138 <= p40_value__138;
    p41_s_0__234 <= p41_s_0__234_comb;
  end

  // ===== Pipe stage 42:
  wire [31:0] p42_temp1__379_comb;
  wire [31:0] p42_e__48_comb;
  wire [12:0] p42_s_1__236_comb;
  wire [9:0] p42_s_1__239_comb;
  wire [6:0] p42_s_1__238_comb;
  wire [1:0] p42_s_1__237_comb;
  wire [5:0] p42_S1__255_comb;
  wire [4:0] p42_S1__254_comb;
  wire [13:0] p42_S1__253_comb;
  wire [6:0] p42_S1__252_comb;
  wire [30:0] p42_add_62492_comb;
  wire [1:0] p42_S0__251_comb;
  wire [10:0] p42_S0__250_comb;
  wire [8:0] p42_S0__249_comb;
  wire [9:0] p42_S0__248_comb;
  wire [31:0] p42_and_62516_comb;
  wire [2:0] p42_s_0__239_comb;
  wire [3:0] p42_s_0__238_comb;
  wire [10:0] p42_s_0__237_comb;
  wire [13:0] p42_s_0__236_comb;
  wire [31:0] p42_S1__48_comb;
  wire [31:0] p42_ch__48_comb;
  wire [31:0] p42_temp1__306_comb;
  wire [31:0] p42_S0__47_comb;
  wire [31:0] p42_maj__47_comb;
  wire [31:0] p42_s_0__240_comb;
  wire [30:0] p42_add_62563_comb;
  wire [31:0] p42_temp1__374_comb;
  wire [31:0] p42_temp1__375_comb;
  wire [31:0] p42_temp2__47_comb;
  wire [30:0] p42_add_62524_comb;
  wire [31:0] p42_temp1__341_comb;
  wire [31:0] p42_temp1__342_comb;
  wire [31:0] p42_temp1__376_comb;
  wire [31:0] p42_a__48_comb;
  wire [31:0] p42_temp1__314_comb;
  wire [31:0] p42_temp1__319_comb;
  wire [31:0] p42_temp1__344_comb;
  assign p42_temp1__379_comb = p41_temp1__377 + p41_temp1__378;
  assign p42_e__48_comb = p41_a__44 + p42_temp1__379_comb;
  assign p42_s_1__236_comb = p41_value__138[29:17] ^ p41_value__138[31:19] ^ p41_value__138[22:10];
  assign p42_s_1__239_comb = p41_value__138[16:7] ^ p41_value__138[18:9];
  assign p42_s_1__238_comb = p41_value__138[6:0] ^ p41_value__138[8:2] ^ p41_value__138[31:25];
  assign p42_s_1__237_comb = p41_value__138[31:30] ^ p41_value__138[1:0] ^ p41_value__138[24:23];
  assign p42_S1__255_comb = p42_e__48_comb[5:0] ^ p42_e__48_comb[10:5] ^ p42_e__48_comb[24:19];
  assign p42_S1__254_comb = p42_e__48_comb[31:27] ^ p42_e__48_comb[4:0] ^ p42_e__48_comb[18:14];
  assign p42_S1__253_comb = p42_e__48_comb[26:13] ^ p42_e__48_comb[31:18] ^ p42_e__48_comb[13:0];
  assign p42_S1__252_comb = p42_e__48_comb[12:6] ^ p42_e__48_comb[17:11] ^ p42_e__48_comb[31:25];
  assign p42_add_62492_comb = p41_value__99[31:1] + 31'h0cd2_608b;
  assign p42_S0__251_comb = p41_a__47[1:0] ^ p41_a__47[12:11] ^ p41_a__47[21:20];
  assign p42_S0__250_comb = p41_a__47[31:21] ^ p41_a__47[10:0] ^ p41_a__47[19:9];
  assign p42_S0__249_comb = p41_a__47[20:12] ^ p41_a__47[31:23] ^ p41_a__47[8:0];
  assign p42_S0__248_comb = p41_a__47[11:2] ^ p41_a__47[22:13] ^ p41_a__47[31:22];
  assign p42_and_62516_comb = p41_a__47 & p41_a__46;
  assign p42_s_0__239_comb = p41_value__99[6:4] ^ p41_value__99[17:15];
  assign p42_s_0__238_comb = p41_value__99[3:0] ^ p41_value__99[14:11] ^ p41_value__99[31:28];
  assign p42_s_0__237_comb = p41_value__99[31:21] ^ p41_value__99[10:0] ^ p41_value__99[27:17];
  assign p42_s_0__236_comb = p41_value__99[20:7] ^ p41_value__99[31:18] ^ p41_value__99[16:3];
  assign p42_S1__48_comb = {p42_S1__255_comb, p42_S1__254_comb, p42_S1__253_comb, p42_S1__252_comb};
  assign p42_ch__48_comb = p42_e__48_comb & p41_e__47 ^ ~(p42_e__48_comb | ~p41_e__46);
  assign p42_temp1__306_comb = {p42_add_62492_comb, p41_value__99[0]};
  assign p42_S0__47_comb = {p42_S0__251_comb, p42_S0__250_comb, p42_S0__249_comb, p42_S0__248_comb};
  assign p42_maj__47_comb = p42_and_62516_comb ^ p41_a__47 & p41_a__45 ^ p41_and_62379;
  assign p42_s_0__240_comb = {p42_s_0__239_comb, p42_s_0__238_comb, p42_s_0__237_comb, p42_s_0__236_comb};
  assign p42_add_62563_comb = {p42_s_1__239_comb, p42_s_1__238_comb, p42_s_1__237_comb, p42_s_1__236_comb[12:1]} + 31'h6338_bc79;
  assign p42_temp1__374_comb = p41_e__45 + p42_S1__48_comb;
  assign p42_temp1__375_comb = p42_ch__48_comb + p42_temp1__306_comb;
  assign p42_temp2__47_comb = p42_S0__47_comb + p42_maj__47_comb;
  assign p42_add_62524_comb = p41_value__123[31:1] + 31'h3a47_c177;
  assign p42_temp1__341_comb = p42_s_0__240_comb + p41_value__123;
  assign p42_temp1__342_comb = {p42_add_62563_comb, p42_s_1__236_comb[0]};
  assign p42_temp1__376_comb = p42_temp1__374_comb + p42_temp1__375_comb;
  assign p42_a__48_comb = p42_temp1__379_comb + p42_temp2__47_comb;
  assign p42_temp1__314_comb = {p42_add_62524_comb, p41_value__123[0]};
  assign p42_temp1__319_comb = p41_value__138 + 32'ha450_6ceb;
  assign p42_temp1__344_comb = p42_temp1__341_comb + p42_temp1__342_comb;

  // Registers for pipe stage 42:
  reg [31:0] p42_e__46;
  reg [31:0] p42_value__93;
  reg [31:0] p42_e__47;
  reg [31:0] p42_value__96;
  reg [31:0] p42_e__48;
  reg [31:0] p42_a__45;
  reg [31:0] p42_temp1__376;
  reg [31:0] p42_temp1__307;
  reg [31:0] p42_a__46;
  reg [31:0] p42_temp1__308;
  reg [31:0] p42_a__47;
  reg [31:0] p42_and_62516;
  reg [31:0] p42_temp1__309;
  reg [31:0] p42_a__48;
  reg [31:0] p42_temp1__310;
  reg [31:0] p42_temp1__311;
  reg [31:0] p42_temp1__312;
  reg [31:0] p42_value__120;
  reg [31:0] p42_temp1__314;
  reg [31:0] p42_temp1__315;
  reg [31:0] p42_temp1__316;
  reg [31:0] p42_temp1__317;
  reg [31:0] p42_value__135;
  reg [31:0] p42_temp1__319;
  reg [3:0] p42_s_0__234;
  reg [31:0] p42_temp1__344;
  always_ff @ (posedge clk) begin
    p42_e__46 <= p41_e__46;
    p42_value__93 <= p41_value__93;
    p42_e__47 <= p41_e__47;
    p42_value__96 <= p41_value__96;
    p42_e__48 <= p42_e__48_comb;
    p42_a__45 <= p41_a__45;
    p42_temp1__376 <= p42_temp1__376_comb;
    p42_temp1__307 <= p41_temp1__307;
    p42_a__46 <= p41_a__46;
    p42_temp1__308 <= p41_temp1__308;
    p42_a__47 <= p41_a__47;
    p42_and_62516 <= p42_and_62516_comb;
    p42_temp1__309 <= p41_temp1__309;
    p42_a__48 <= p42_a__48_comb;
    p42_temp1__310 <= p41_temp1__310;
    p42_temp1__311 <= p41_temp1__311;
    p42_temp1__312 <= p41_temp1__312;
    p42_value__120 <= p41_value__120;
    p42_temp1__314 <= p42_temp1__314_comb;
    p42_temp1__315 <= p41_temp1__315;
    p42_temp1__316 <= p41_temp1__316;
    p42_temp1__317 <= p41_temp1__317;
    p42_value__135 <= p41_value__135;
    p42_temp1__319 <= p42_temp1__319_comb;
    p42_s_0__234 <= p41_s_0__234;
    p42_temp1__344 <= p42_temp1__344_comb;
  end

  // ===== Pipe stage 43:
  wire [1:0] p43_S0__255_comb;
  wire [10:0] p43_S0__254_comb;
  wire [8:0] p43_S0__253_comb;
  wire [9:0] p43_S0__252_comb;
  wire [31:0] p43_and_62662_comb;
  wire [31:0] p43_S0__48_comb;
  wire [31:0] p43_maj__48_comb;
  wire [31:0] p43_e__49_comb;
  wire [31:0] p43_temp2__48_comb;
  wire [31:0] p43_a__49_comb;
  wire [5:0] p43_S1__259_comb;
  wire [4:0] p43_S1__258_comb;
  wire [13:0] p43_S1__257_comb;
  wire [6:0] p43_S1__256_comb;
  wire [31:0] p43_S1__49_comb;
  wire [31:0] p43_ch__49_comb;
  wire [1:0] p43_S0__259_comb;
  wire [10:0] p43_S0__258_comb;
  wire [8:0] p43_S0__257_comb;
  wire [9:0] p43_S0__256_comb;
  wire [31:0] p43_and_62684_comb;
  wire [31:0] p43_temp1__371_comb;
  wire [31:0] p43_temp1__372_comb;
  wire [31:0] p43_S0__49_comb;
  wire [31:0] p43_maj__49_comb;
  wire [31:0] p43_temp1__373_comb;
  wire [31:0] p43_temp2__49_comb;
  wire [31:0] p43_e__50_comb;
  wire [31:0] p43_a__50_comb;
  assign p43_S0__255_comb = p42_a__48[1:0] ^ p42_a__48[12:11] ^ p42_a__48[21:20];
  assign p43_S0__254_comb = p42_a__48[31:21] ^ p42_a__48[10:0] ^ p42_a__48[19:9];
  assign p43_S0__253_comb = p42_a__48[20:12] ^ p42_a__48[31:23] ^ p42_a__48[8:0];
  assign p43_S0__252_comb = p42_a__48[11:2] ^ p42_a__48[22:13] ^ p42_a__48[31:22];
  assign p43_and_62662_comb = p42_a__48 & p42_a__47;
  assign p43_S0__48_comb = {p43_S0__255_comb, p43_S0__254_comb, p43_S0__253_comb, p43_S0__252_comb};
  assign p43_maj__48_comb = p43_and_62662_comb ^ p42_a__48 & p42_a__46 ^ p42_and_62516;
  assign p43_e__49_comb = p42_a__45 + p42_temp1__376;
  assign p43_temp2__48_comb = p43_S0__48_comb + p43_maj__48_comb;
  assign p43_a__49_comb = p42_temp1__376 + p43_temp2__48_comb;
  assign p43_S1__259_comb = p43_e__49_comb[5:0] ^ p43_e__49_comb[10:5] ^ p43_e__49_comb[24:19];
  assign p43_S1__258_comb = p43_e__49_comb[31:27] ^ p43_e__49_comb[4:0] ^ p43_e__49_comb[18:14];
  assign p43_S1__257_comb = p43_e__49_comb[26:13] ^ p43_e__49_comb[31:18] ^ p43_e__49_comb[13:0];
  assign p43_S1__256_comb = p43_e__49_comb[12:6] ^ p43_e__49_comb[17:11] ^ p43_e__49_comb[31:25];
  assign p43_S1__49_comb = {p43_S1__259_comb, p43_S1__258_comb, p43_S1__257_comb, p43_S1__256_comb};
  assign p43_ch__49_comb = p43_e__49_comb & p42_e__48 ^ ~(p43_e__49_comb | ~p42_e__47);
  assign p43_S0__259_comb = p43_a__49_comb[1:0] ^ p43_a__49_comb[12:11] ^ p43_a__49_comb[21:20];
  assign p43_S0__258_comb = p43_a__49_comb[31:21] ^ p43_a__49_comb[10:0] ^ p43_a__49_comb[19:9];
  assign p43_S0__257_comb = p43_a__49_comb[20:12] ^ p43_a__49_comb[31:23] ^ p43_a__49_comb[8:0];
  assign p43_S0__256_comb = p43_a__49_comb[11:2] ^ p43_a__49_comb[22:13] ^ p43_a__49_comb[31:22];
  assign p43_and_62684_comb = p43_a__49_comb & p42_a__48;
  assign p43_temp1__371_comb = p42_e__46 + p43_S1__49_comb;
  assign p43_temp1__372_comb = p43_ch__49_comb + p42_temp1__307;
  assign p43_S0__49_comb = {p43_S0__259_comb, p43_S0__258_comb, p43_S0__257_comb, p43_S0__256_comb};
  assign p43_maj__49_comb = p43_and_62684_comb ^ p43_a__49_comb & p42_a__47 ^ p43_and_62662_comb;
  assign p43_temp1__373_comb = p43_temp1__371_comb + p43_temp1__372_comb;
  assign p43_temp2__49_comb = p43_S0__49_comb + p43_maj__49_comb;
  assign p43_e__50_comb = p42_a__46 + p43_temp1__373_comb;
  assign p43_a__50_comb = p43_temp1__373_comb + p43_temp2__49_comb;

  // Registers for pipe stage 43:
  reg [31:0] p43_value__93;
  reg [31:0] p43_e__47;
  reg [31:0] p43_value__96;
  reg [31:0] p43_e__48;
  reg [31:0] p43_e__49;
  reg [31:0] p43_e__50;
  reg [31:0] p43_temp1__308;
  reg [31:0] p43_a__47;
  reg [31:0] p43_temp1__309;
  reg [31:0] p43_a__48;
  reg [31:0] p43_temp1__310;
  reg [31:0] p43_a__49;
  reg [31:0] p43_and_62684;
  reg [31:0] p43_temp1__311;
  reg [31:0] p43_a__50;
  reg [31:0] p43_temp1__312;
  reg [31:0] p43_value__120;
  reg [31:0] p43_temp1__314;
  reg [31:0] p43_temp1__315;
  reg [31:0] p43_temp1__316;
  reg [31:0] p43_temp1__317;
  reg [31:0] p43_value__135;
  reg [31:0] p43_temp1__319;
  reg [3:0] p43_s_0__234;
  reg [31:0] p43_temp1__344;
  always_ff @ (posedge clk) begin
    p43_value__93 <= p42_value__93;
    p43_e__47 <= p42_e__47;
    p43_value__96 <= p42_value__96;
    p43_e__48 <= p42_e__48;
    p43_e__49 <= p43_e__49_comb;
    p43_e__50 <= p43_e__50_comb;
    p43_temp1__308 <= p42_temp1__308;
    p43_a__47 <= p42_a__47;
    p43_temp1__309 <= p42_temp1__309;
    p43_a__48 <= p42_a__48;
    p43_temp1__310 <= p42_temp1__310;
    p43_a__49 <= p43_a__49_comb;
    p43_and_62684 <= p43_and_62684_comb;
    p43_temp1__311 <= p42_temp1__311;
    p43_a__50 <= p43_a__50_comb;
    p43_temp1__312 <= p42_temp1__312;
    p43_value__120 <= p42_value__120;
    p43_temp1__314 <= p42_temp1__314;
    p43_temp1__315 <= p42_temp1__315;
    p43_temp1__316 <= p42_temp1__316;
    p43_temp1__317 <= p42_temp1__317;
    p43_value__135 <= p42_value__135;
    p43_temp1__319 <= p42_temp1__319;
    p43_s_0__234 <= p42_s_0__234;
    p43_temp1__344 <= p42_temp1__344;
  end

  // ===== Pipe stage 44:
  wire [5:0] p44_S1__263_comb;
  wire [4:0] p44_S1__262_comb;
  wire [13:0] p44_S1__261_comb;
  wire [6:0] p44_S1__260_comb;
  wire [31:0] p44_S1__50_comb;
  wire [31:0] p44_ch__50_comb;
  wire [31:0] p44_temp1__368_comb;
  wire [31:0] p44_temp1__369_comb;
  wire [31:0] p44_temp1__370_comb;
  wire [31:0] p44_e__51_comb;
  wire [1:0] p44_S0__263_comb;
  wire [10:0] p44_S0__262_comb;
  wire [8:0] p44_S0__261_comb;
  wire [9:0] p44_S0__260_comb;
  wire [31:0] p44_and_62799_comb;
  wire [5:0] p44_S1__267_comb;
  wire [4:0] p44_S1__266_comb;
  wire [13:0] p44_S1__265_comb;
  wire [6:0] p44_S1__264_comb;
  wire [31:0] p44_S0__50_comb;
  wire [31:0] p44_maj__50_comb;
  wire [31:0] p44_S1__51_comb;
  wire [31:0] p44_temp2__50_comb;
  wire [31:0] p44_temp1__205_comb;
  wire [31:0] p44_a__51_comb;
  assign p44_S1__263_comb = p43_e__50[5:0] ^ p43_e__50[10:5] ^ p43_e__50[24:19];
  assign p44_S1__262_comb = p43_e__50[31:27] ^ p43_e__50[4:0] ^ p43_e__50[18:14];
  assign p44_S1__261_comb = p43_e__50[26:13] ^ p43_e__50[31:18] ^ p43_e__50[13:0];
  assign p44_S1__260_comb = p43_e__50[12:6] ^ p43_e__50[17:11] ^ p43_e__50[31:25];
  assign p44_S1__50_comb = {p44_S1__263_comb, p44_S1__262_comb, p44_S1__261_comb, p44_S1__260_comb};
  assign p44_ch__50_comb = p43_e__50 & p43_e__49 ^ ~(p43_e__50 | ~p43_e__48);
  assign p44_temp1__368_comb = p43_e__47 + p44_S1__50_comb;
  assign p44_temp1__369_comb = p44_ch__50_comb + p43_temp1__308;
  assign p44_temp1__370_comb = p44_temp1__368_comb + p44_temp1__369_comb;
  assign p44_e__51_comb = p43_a__47 + p44_temp1__370_comb;
  assign p44_S0__263_comb = p43_a__50[1:0] ^ p43_a__50[12:11] ^ p43_a__50[21:20];
  assign p44_S0__262_comb = p43_a__50[31:21] ^ p43_a__50[10:0] ^ p43_a__50[19:9];
  assign p44_S0__261_comb = p43_a__50[20:12] ^ p43_a__50[31:23] ^ p43_a__50[8:0];
  assign p44_S0__260_comb = p43_a__50[11:2] ^ p43_a__50[22:13] ^ p43_a__50[31:22];
  assign p44_and_62799_comb = p43_a__50 & p43_a__49;
  assign p44_S1__267_comb = p44_e__51_comb[5:0] ^ p44_e__51_comb[10:5] ^ p44_e__51_comb[24:19];
  assign p44_S1__266_comb = p44_e__51_comb[31:27] ^ p44_e__51_comb[4:0] ^ p44_e__51_comb[18:14];
  assign p44_S1__265_comb = p44_e__51_comb[26:13] ^ p44_e__51_comb[31:18] ^ p44_e__51_comb[13:0];
  assign p44_S1__264_comb = p44_e__51_comb[12:6] ^ p44_e__51_comb[17:11] ^ p44_e__51_comb[31:25];
  assign p44_S0__50_comb = {p44_S0__263_comb, p44_S0__262_comb, p44_S0__261_comb, p44_S0__260_comb};
  assign p44_maj__50_comb = p44_and_62799_comb ^ p43_a__50 & p43_a__48 ^ p43_and_62684;
  assign p44_S1__51_comb = {p44_S1__267_comb, p44_S1__266_comb, p44_S1__265_comb, p44_S1__264_comb};
  assign p44_temp2__50_comb = p44_S0__50_comb + p44_maj__50_comb;
  assign p44_temp1__205_comb = p43_e__48 + p44_S1__51_comb;
  assign p44_a__51_comb = p44_temp1__370_comb + p44_temp2__50_comb;

  // Registers for pipe stage 44:
  reg [31:0] p44_value__93;
  reg [31:0] p44_value__96;
  reg [31:0] p44_e__49;
  reg [31:0] p44_e__50;
  reg [31:0] p44_e__51;
  reg [31:0] p44_temp1__205;
  reg [31:0] p44_temp1__309;
  reg [31:0] p44_a__48;
  reg [31:0] p44_temp1__310;
  reg [31:0] p44_a__49;
  reg [31:0] p44_temp1__311;
  reg [31:0] p44_a__50;
  reg [31:0] p44_and_62799;
  reg [31:0] p44_a__51;
  reg [31:0] p44_temp1__312;
  reg [31:0] p44_value__120;
  reg [31:0] p44_temp1__314;
  reg [31:0] p44_temp1__315;
  reg [31:0] p44_temp1__316;
  reg [31:0] p44_temp1__317;
  reg [31:0] p44_value__135;
  reg [31:0] p44_temp1__319;
  reg [3:0] p44_s_0__234;
  reg [31:0] p44_temp1__344;
  always_ff @ (posedge clk) begin
    p44_value__93 <= p43_value__93;
    p44_value__96 <= p43_value__96;
    p44_e__49 <= p43_e__49;
    p44_e__50 <= p43_e__50;
    p44_e__51 <= p44_e__51_comb;
    p44_temp1__205 <= p44_temp1__205_comb;
    p44_temp1__309 <= p43_temp1__309;
    p44_a__48 <= p43_a__48;
    p44_temp1__310 <= p43_temp1__310;
    p44_a__49 <= p43_a__49;
    p44_temp1__311 <= p43_temp1__311;
    p44_a__50 <= p43_a__50;
    p44_and_62799 <= p44_and_62799_comb;
    p44_a__51 <= p44_a__51_comb;
    p44_temp1__312 <= p43_temp1__312;
    p44_value__120 <= p43_value__120;
    p44_temp1__314 <= p43_temp1__314;
    p44_temp1__315 <= p43_temp1__315;
    p44_temp1__316 <= p43_temp1__316;
    p44_temp1__317 <= p43_temp1__317;
    p44_value__135 <= p43_value__135;
    p44_temp1__319 <= p43_temp1__319;
    p44_s_0__234 <= p43_s_0__234;
    p44_temp1__344 <= p43_temp1__344;
  end

  // ===== Pipe stage 45:
  wire [31:0] p45_ch__51_comb;
  wire [31:0] p45_temp1__206_comb;
  wire [31:0] p45_temp1__208_comb;
  wire [31:0] p45_e__52_comb;
  wire [1:0] p45_S0__267_comb;
  wire [10:0] p45_S0__266_comb;
  wire [8:0] p45_S0__265_comb;
  wire [9:0] p45_S0__264_comb;
  wire [31:0] p45_and_62894_comb;
  wire [5:0] p45_S1__271_comb;
  wire [4:0] p45_S1__270_comb;
  wire [13:0] p45_S1__269_comb;
  wire [6:0] p45_S1__268_comb;
  wire [31:0] p45_S0__51_comb;
  wire [31:0] p45_maj__51_comb;
  wire [31:0] p45_S1__52_comb;
  wire [31:0] p45_temp2__51_comb;
  wire [31:0] p45_temp1__209_comb;
  wire [31:0] p45_a__52_comb;
  assign p45_ch__51_comb = p44_e__51 & p44_e__50 ^ ~(p44_e__51 | ~p44_e__49);
  assign p45_temp1__206_comb = p44_temp1__205 + p45_ch__51_comb;
  assign p45_temp1__208_comb = p45_temp1__206_comb + p44_temp1__309;
  assign p45_e__52_comb = p44_a__48 + p45_temp1__208_comb;
  assign p45_S0__267_comb = p44_a__51[1:0] ^ p44_a__51[12:11] ^ p44_a__51[21:20];
  assign p45_S0__266_comb = p44_a__51[31:21] ^ p44_a__51[10:0] ^ p44_a__51[19:9];
  assign p45_S0__265_comb = p44_a__51[20:12] ^ p44_a__51[31:23] ^ p44_a__51[8:0];
  assign p45_S0__264_comb = p44_a__51[11:2] ^ p44_a__51[22:13] ^ p44_a__51[31:22];
  assign p45_and_62894_comb = p44_a__51 & p44_a__50;
  assign p45_S1__271_comb = p45_e__52_comb[5:0] ^ p45_e__52_comb[10:5] ^ p45_e__52_comb[24:19];
  assign p45_S1__270_comb = p45_e__52_comb[31:27] ^ p45_e__52_comb[4:0] ^ p45_e__52_comb[18:14];
  assign p45_S1__269_comb = p45_e__52_comb[26:13] ^ p45_e__52_comb[31:18] ^ p45_e__52_comb[13:0];
  assign p45_S1__268_comb = p45_e__52_comb[12:6] ^ p45_e__52_comb[17:11] ^ p45_e__52_comb[31:25];
  assign p45_S0__51_comb = {p45_S0__267_comb, p45_S0__266_comb, p45_S0__265_comb, p45_S0__264_comb};
  assign p45_maj__51_comb = p45_and_62894_comb ^ p44_a__51 & p44_a__49 ^ p44_and_62799;
  assign p45_S1__52_comb = {p45_S1__271_comb, p45_S1__270_comb, p45_S1__269_comb, p45_S1__268_comb};
  assign p45_temp2__51_comb = p45_S0__51_comb + p45_maj__51_comb;
  assign p45_temp1__209_comb = p44_e__49 + p45_S1__52_comb;
  assign p45_a__52_comb = p45_temp1__208_comb + p45_temp2__51_comb;

  // Registers for pipe stage 45:
  reg [31:0] p45_value__93;
  reg [31:0] p45_value__96;
  reg [31:0] p45_e__50;
  reg [31:0] p45_e__51;
  reg [31:0] p45_e__52;
  reg [31:0] p45_temp1__209;
  reg [31:0] p45_temp1__310;
  reg [31:0] p45_a__49;
  reg [31:0] p45_temp1__311;
  reg [31:0] p45_a__50;
  reg [31:0] p45_a__51;
  reg [31:0] p45_and_62894;
  reg [31:0] p45_temp1__312;
  reg [31:0] p45_a__52;
  reg [31:0] p45_value__120;
  reg [31:0] p45_temp1__314;
  reg [31:0] p45_temp1__315;
  reg [31:0] p45_temp1__316;
  reg [31:0] p45_temp1__317;
  reg [31:0] p45_value__135;
  reg [31:0] p45_temp1__319;
  reg [3:0] p45_s_0__234;
  reg [31:0] p45_temp1__344;
  always_ff @ (posedge clk) begin
    p45_value__93 <= p44_value__93;
    p45_value__96 <= p44_value__96;
    p45_e__50 <= p44_e__50;
    p45_e__51 <= p44_e__51;
    p45_e__52 <= p45_e__52_comb;
    p45_temp1__209 <= p45_temp1__209_comb;
    p45_temp1__310 <= p44_temp1__310;
    p45_a__49 <= p44_a__49;
    p45_temp1__311 <= p44_temp1__311;
    p45_a__50 <= p44_a__50;
    p45_a__51 <= p44_a__51;
    p45_and_62894 <= p45_and_62894_comb;
    p45_temp1__312 <= p44_temp1__312;
    p45_a__52 <= p45_a__52_comb;
    p45_value__120 <= p44_value__120;
    p45_temp1__314 <= p44_temp1__314;
    p45_temp1__315 <= p44_temp1__315;
    p45_temp1__316 <= p44_temp1__316;
    p45_temp1__317 <= p44_temp1__317;
    p45_value__135 <= p44_value__135;
    p45_temp1__319 <= p44_temp1__319;
    p45_s_0__234 <= p44_s_0__234;
    p45_temp1__344 <= p44_temp1__344;
  end

  // ===== Pipe stage 46:
  wire [31:0] p46_ch__52_comb;
  wire [31:0] p46_temp1__210_comb;
  wire [31:0] p46_temp1__212_comb;
  wire [31:0] p46_e__53_comb;
  wire [1:0] p46_S0__271_comb;
  wire [10:0] p46_S0__270_comb;
  wire [8:0] p46_S0__269_comb;
  wire [9:0] p46_S0__268_comb;
  wire [31:0] p46_and_62992_comb;
  wire [5:0] p46_S1__275_comb;
  wire [4:0] p46_S1__274_comb;
  wire [13:0] p46_S1__273_comb;
  wire [6:0] p46_S1__272_comb;
  wire [31:0] p46_S0__52_comb;
  wire [31:0] p46_maj__52_comb;
  wire [31:0] p46_S1__53_comb;
  wire [31:0] p46_ch__53_comb;
  wire [31:0] p46_temp2__52_comb;
  wire [31:0] p46_temp1__365_comb;
  wire [31:0] p46_temp1__366_comb;
  wire [31:0] p46_a__53_comb;
  assign p46_ch__52_comb = p45_e__52 & p45_e__51 ^ ~(p45_e__52 | ~p45_e__50);
  assign p46_temp1__210_comb = p45_temp1__209 + p46_ch__52_comb;
  assign p46_temp1__212_comb = p46_temp1__210_comb + p45_temp1__310;
  assign p46_e__53_comb = p45_a__49 + p46_temp1__212_comb;
  assign p46_S0__271_comb = p45_a__52[1:0] ^ p45_a__52[12:11] ^ p45_a__52[21:20];
  assign p46_S0__270_comb = p45_a__52[31:21] ^ p45_a__52[10:0] ^ p45_a__52[19:9];
  assign p46_S0__269_comb = p45_a__52[20:12] ^ p45_a__52[31:23] ^ p45_a__52[8:0];
  assign p46_S0__268_comb = p45_a__52[11:2] ^ p45_a__52[22:13] ^ p45_a__52[31:22];
  assign p46_and_62992_comb = p45_a__52 & p45_a__51;
  assign p46_S1__275_comb = p46_e__53_comb[5:0] ^ p46_e__53_comb[10:5] ^ p46_e__53_comb[24:19];
  assign p46_S1__274_comb = p46_e__53_comb[31:27] ^ p46_e__53_comb[4:0] ^ p46_e__53_comb[18:14];
  assign p46_S1__273_comb = p46_e__53_comb[26:13] ^ p46_e__53_comb[31:18] ^ p46_e__53_comb[13:0];
  assign p46_S1__272_comb = p46_e__53_comb[12:6] ^ p46_e__53_comb[17:11] ^ p46_e__53_comb[31:25];
  assign p46_S0__52_comb = {p46_S0__271_comb, p46_S0__270_comb, p46_S0__269_comb, p46_S0__268_comb};
  assign p46_maj__52_comb = p46_and_62992_comb ^ p45_a__52 & p45_a__50 ^ p45_and_62894;
  assign p46_S1__53_comb = {p46_S1__275_comb, p46_S1__274_comb, p46_S1__273_comb, p46_S1__272_comb};
  assign p46_ch__53_comb = p46_e__53_comb & p45_e__52 ^ ~(p46_e__53_comb | ~p45_e__51);
  assign p46_temp2__52_comb = p46_S0__52_comb + p46_maj__52_comb;
  assign p46_temp1__365_comb = p45_e__50 + p46_S1__53_comb;
  assign p46_temp1__366_comb = p46_ch__53_comb + p45_temp1__311;
  assign p46_a__53_comb = p46_temp1__212_comb + p46_temp2__52_comb;

  // Registers for pipe stage 46:
  reg [31:0] p46_value__93;
  reg [31:0] p46_value__96;
  reg [31:0] p46_e__51;
  reg [31:0] p46_e__52;
  reg [31:0] p46_e__53;
  reg [31:0] p46_a__50;
  reg [31:0] p46_temp1__365;
  reg [31:0] p46_temp1__366;
  reg [31:0] p46_a__51;
  reg [31:0] p46_temp1__312;
  reg [31:0] p46_a__52;
  reg [31:0] p46_and_62992;
  reg [31:0] p46_value__120;
  reg [31:0] p46_a__53;
  reg [31:0] p46_temp1__314;
  reg [31:0] p46_temp1__315;
  reg [31:0] p46_temp1__316;
  reg [31:0] p46_temp1__317;
  reg [31:0] p46_value__135;
  reg [31:0] p46_temp1__319;
  reg [3:0] p46_s_0__234;
  reg [31:0] p46_temp1__344;
  always_ff @ (posedge clk) begin
    p46_value__93 <= p45_value__93;
    p46_value__96 <= p45_value__96;
    p46_e__51 <= p45_e__51;
    p46_e__52 <= p45_e__52;
    p46_e__53 <= p46_e__53_comb;
    p46_a__50 <= p45_a__50;
    p46_temp1__365 <= p46_temp1__365_comb;
    p46_temp1__366 <= p46_temp1__366_comb;
    p46_a__51 <= p45_a__51;
    p46_temp1__312 <= p45_temp1__312;
    p46_a__52 <= p45_a__52;
    p46_and_62992 <= p46_and_62992_comb;
    p46_value__120 <= p45_value__120;
    p46_a__53 <= p46_a__53_comb;
    p46_temp1__314 <= p45_temp1__314;
    p46_temp1__315 <= p45_temp1__315;
    p46_temp1__316 <= p45_temp1__316;
    p46_temp1__317 <= p45_temp1__317;
    p46_value__135 <= p45_value__135;
    p46_temp1__319 <= p45_temp1__319;
    p46_s_0__234 <= p45_s_0__234;
    p46_temp1__344 <= p45_temp1__344;
  end

  // ===== Pipe stage 47:
  wire [31:0] p47_temp1__367_comb;
  wire [31:0] p47_e__54_comb;
  wire [5:0] p47_S1__279_comb;
  wire [4:0] p47_S1__278_comb;
  wire [13:0] p47_S1__277_comb;
  wire [6:0] p47_S1__276_comb;
  wire [1:0] p47_S0__275_comb;
  wire [10:0] p47_S0__274_comb;
  wire [8:0] p47_S0__273_comb;
  wire [9:0] p47_S0__272_comb;
  wire [31:0] p47_and_63083_comb;
  wire [31:0] p47_S1__54_comb;
  wire [31:0] p47_S0__53_comb;
  wire [31:0] p47_maj__53_comb;
  wire [31:0] p47_temp1__217_comb;
  wire [31:0] p47_ch__54_comb;
  wire [31:0] p47_temp2__53_comb;
  wire [31:0] p47_temp1__218_comb;
  wire [31:0] p47_a__54_comb;
  assign p47_temp1__367_comb = p46_temp1__365 + p46_temp1__366;
  assign p47_e__54_comb = p46_a__50 + p47_temp1__367_comb;
  assign p47_S1__279_comb = p47_e__54_comb[5:0] ^ p47_e__54_comb[10:5] ^ p47_e__54_comb[24:19];
  assign p47_S1__278_comb = p47_e__54_comb[31:27] ^ p47_e__54_comb[4:0] ^ p47_e__54_comb[18:14];
  assign p47_S1__277_comb = p47_e__54_comb[26:13] ^ p47_e__54_comb[31:18] ^ p47_e__54_comb[13:0];
  assign p47_S1__276_comb = p47_e__54_comb[12:6] ^ p47_e__54_comb[17:11] ^ p47_e__54_comb[31:25];
  assign p47_S0__275_comb = p46_a__53[1:0] ^ p46_a__53[12:11] ^ p46_a__53[21:20];
  assign p47_S0__274_comb = p46_a__53[31:21] ^ p46_a__53[10:0] ^ p46_a__53[19:9];
  assign p47_S0__273_comb = p46_a__53[20:12] ^ p46_a__53[31:23] ^ p46_a__53[8:0];
  assign p47_S0__272_comb = p46_a__53[11:2] ^ p46_a__53[22:13] ^ p46_a__53[31:22];
  assign p47_and_63083_comb = p46_a__53 & p46_a__52;
  assign p47_S1__54_comb = {p47_S1__279_comb, p47_S1__278_comb, p47_S1__277_comb, p47_S1__276_comb};
  assign p47_S0__53_comb = {p47_S0__275_comb, p47_S0__274_comb, p47_S0__273_comb, p47_S0__272_comb};
  assign p47_maj__53_comb = p47_and_63083_comb ^ p46_a__53 & p46_a__51 ^ p46_and_62992;
  assign p47_temp1__217_comb = p46_e__51 + p47_S1__54_comb;
  assign p47_ch__54_comb = p47_e__54_comb & p46_e__53 ^ ~(p47_e__54_comb | ~p46_e__52);
  assign p47_temp2__53_comb = p47_S0__53_comb + p47_maj__53_comb;
  assign p47_temp1__218_comb = p47_temp1__217_comb + p47_ch__54_comb;
  assign p47_a__54_comb = p47_temp1__367_comb + p47_temp2__53_comb;

  // Registers for pipe stage 47:
  reg [31:0] p47_value__93;
  reg [31:0] p47_value__96;
  reg [31:0] p47_e__52;
  reg [31:0] p47_e__53;
  reg [31:0] p47_e__54;
  reg [31:0] p47_a__51;
  reg [31:0] p47_temp1__218;
  reg [31:0] p47_temp1__312;
  reg [31:0] p47_a__52;
  reg [31:0] p47_value__120;
  reg [31:0] p47_a__53;
  reg [31:0] p47_and_63083;
  reg [31:0] p47_temp1__314;
  reg [31:0] p47_a__54;
  reg [31:0] p47_temp1__315;
  reg [31:0] p47_temp1__316;
  reg [31:0] p47_temp1__317;
  reg [31:0] p47_value__135;
  reg [31:0] p47_temp1__319;
  reg [3:0] p47_s_0__234;
  reg [31:0] p47_temp1__344;
  always_ff @ (posedge clk) begin
    p47_value__93 <= p46_value__93;
    p47_value__96 <= p46_value__96;
    p47_e__52 <= p46_e__52;
    p47_e__53 <= p46_e__53;
    p47_e__54 <= p47_e__54_comb;
    p47_a__51 <= p46_a__51;
    p47_temp1__218 <= p47_temp1__218_comb;
    p47_temp1__312 <= p46_temp1__312;
    p47_a__52 <= p46_a__52;
    p47_value__120 <= p46_value__120;
    p47_a__53 <= p46_a__53;
    p47_and_63083 <= p47_and_63083_comb;
    p47_temp1__314 <= p46_temp1__314;
    p47_a__54 <= p47_a__54_comb;
    p47_temp1__315 <= p46_temp1__315;
    p47_temp1__316 <= p46_temp1__316;
    p47_temp1__317 <= p46_temp1__317;
    p47_value__135 <= p46_value__135;
    p47_temp1__319 <= p46_temp1__319;
    p47_s_0__234 <= p46_s_0__234;
    p47_temp1__344 <= p46_temp1__344;
  end

  // ===== Pipe stage 48:
  wire [31:0] p48_temp1__220_comb;
  wire [31:0] p48_e__55_comb;
  wire [5:0] p48_S1__283_comb;
  wire [4:0] p48_S1__282_comb;
  wire [13:0] p48_S1__281_comb;
  wire [6:0] p48_S1__280_comb;
  wire [1:0] p48_S0__279_comb;
  wire [10:0] p48_S0__278_comb;
  wire [8:0] p48_S0__277_comb;
  wire [9:0] p48_S0__276_comb;
  wire [31:0] p48_and_63174_comb;
  wire [2:0] p48_s_0__235_comb;
  wire [10:0] p48_s_0__233_comb;
  wire [13:0] p48_s_0__232_comb;
  wire [9:0] p48_s_1__235_comb;
  wire [6:0] p48_s_1__234_comb;
  wire [1:0] p48_s_1__233_comb;
  wire [12:0] p48_s_1__232_comb;
  wire [31:0] p48_S1__55_comb;
  wire [31:0] p48_S0__54_comb;
  wire [31:0] p48_maj__54_comb;
  wire [31:0] p48_s_0__47_comb;
  wire [31:0] p48_s_1__47_comb;
  wire [31:0] p48_temp1__221_comb;
  wire [31:0] p48_ch__55_comb;
  wire [31:0] p48_temp2__54_comb;
  wire [30:0] p48_add_63182_comb;
  wire [31:0] p48_temp1__348_comb;
  wire [31:0] p48_temp1__349_comb;
  wire [31:0] p48_temp1__222_comb;
  wire [31:0] p48_temp1__313_comb;
  wire [31:0] p48_a__55_comb;
  wire [31:0] p48_temp1__318_comb;
  wire [31:0] p48_temp1__351_comb;
  assign p48_temp1__220_comb = p47_temp1__218 + p47_temp1__312;
  assign p48_e__55_comb = p47_a__51 + p48_temp1__220_comb;
  assign p48_S1__283_comb = p48_e__55_comb[5:0] ^ p48_e__55_comb[10:5] ^ p48_e__55_comb[24:19];
  assign p48_S1__282_comb = p48_e__55_comb[31:27] ^ p48_e__55_comb[4:0] ^ p48_e__55_comb[18:14];
  assign p48_S1__281_comb = p48_e__55_comb[26:13] ^ p48_e__55_comb[31:18] ^ p48_e__55_comb[13:0];
  assign p48_S1__280_comb = p48_e__55_comb[12:6] ^ p48_e__55_comb[17:11] ^ p48_e__55_comb[31:25];
  assign p48_S0__279_comb = p47_a__54[1:0] ^ p47_a__54[12:11] ^ p47_a__54[21:20];
  assign p48_S0__278_comb = p47_a__54[31:21] ^ p47_a__54[10:0] ^ p47_a__54[19:9];
  assign p48_S0__277_comb = p47_a__54[20:12] ^ p47_a__54[31:23] ^ p47_a__54[8:0];
  assign p48_S0__276_comb = p47_a__54[11:2] ^ p47_a__54[22:13] ^ p47_a__54[31:22];
  assign p48_and_63174_comb = p47_a__54 & p47_a__53;
  assign p48_s_0__235_comb = p47_value__96[6:4] ^ p47_value__96[17:15];
  assign p48_s_0__233_comb = p47_value__96[31:21] ^ p47_value__96[10:0] ^ p47_value__96[27:17];
  assign p48_s_0__232_comb = p47_value__96[20:7] ^ p47_value__96[31:18] ^ p47_value__96[16:3];
  assign p48_s_1__235_comb = p47_value__135[16:7] ^ p47_value__135[18:9];
  assign p48_s_1__234_comb = p47_value__135[6:0] ^ p47_value__135[8:2] ^ p47_value__135[31:25];
  assign p48_s_1__233_comb = p47_value__135[31:30] ^ p47_value__135[1:0] ^ p47_value__135[24:23];
  assign p48_s_1__232_comb = p47_value__135[29:17] ^ p47_value__135[31:19] ^ p47_value__135[22:10];
  assign p48_S1__55_comb = {p48_S1__283_comb, p48_S1__282_comb, p48_S1__281_comb, p48_S1__280_comb};
  assign p48_S0__54_comb = {p48_S0__279_comb, p48_S0__278_comb, p48_S0__277_comb, p48_S0__276_comb};
  assign p48_maj__54_comb = p48_and_63174_comb ^ p47_a__54 & p47_a__52 ^ p47_and_63083;
  assign p48_s_0__47_comb = {p48_s_0__235_comb, p47_s_0__234, p48_s_0__233_comb, p48_s_0__232_comb};
  assign p48_s_1__47_comb = {p48_s_1__235_comb, p48_s_1__234_comb, p48_s_1__233_comb, p48_s_1__232_comb};
  assign p48_temp1__221_comb = p47_e__52 + p48_S1__55_comb;
  assign p48_ch__55_comb = p48_e__55_comb & p47_e__54 ^ ~(p48_e__55_comb | ~p47_e__53);
  assign p48_temp2__54_comb = p48_S0__54_comb + p48_maj__54_comb;
  assign p48_add_63182_comb = p47_value__135[31:1] + 31'h485f_7ffd;
  assign p48_temp1__348_comb = p48_s_0__47_comb + p47_value__120;
  assign p48_temp1__349_comb = p48_s_1__47_comb + 32'hbef9_a3f7;
  assign p48_temp1__222_comb = p48_temp1__221_comb + p48_ch__55_comb;
  assign p48_temp1__313_comb = p47_value__120 + 32'h682e_6ff3;
  assign p48_a__55_comb = p48_temp1__220_comb + p48_temp2__54_comb;
  assign p48_temp1__318_comb = {p48_add_63182_comb, p47_value__135[0]};
  assign p48_temp1__351_comb = p48_temp1__348_comb + p48_temp1__349_comb;

  // Registers for pipe stage 48:
  reg [31:0] p48_value__93;
  reg [31:0] p48_value__96;
  reg [31:0] p48_e__53;
  reg [31:0] p48_e__54;
  reg [31:0] p48_e__55;
  reg [31:0] p48_a__52;
  reg [31:0] p48_temp1__222;
  reg [31:0] p48_temp1__313;
  reg [31:0] p48_a__53;
  reg [31:0] p48_temp1__314;
  reg [31:0] p48_a__54;
  reg [31:0] p48_and_63174;
  reg [31:0] p48_a__55;
  reg [31:0] p48_temp1__315;
  reg [31:0] p48_temp1__316;
  reg [31:0] p48_temp1__317;
  reg [31:0] p48_temp1__318;
  reg [31:0] p48_temp1__319;
  reg [31:0] p48_temp1__351;
  reg [31:0] p48_temp1__344;
  always_ff @ (posedge clk) begin
    p48_value__93 <= p47_value__93;
    p48_value__96 <= p47_value__96;
    p48_e__53 <= p47_e__53;
    p48_e__54 <= p47_e__54;
    p48_e__55 <= p48_e__55_comb;
    p48_a__52 <= p47_a__52;
    p48_temp1__222 <= p48_temp1__222_comb;
    p48_temp1__313 <= p48_temp1__313_comb;
    p48_a__53 <= p47_a__53;
    p48_temp1__314 <= p47_temp1__314;
    p48_a__54 <= p47_a__54;
    p48_and_63174 <= p48_and_63174_comb;
    p48_a__55 <= p48_a__55_comb;
    p48_temp1__315 <= p47_temp1__315;
    p48_temp1__316 <= p47_temp1__316;
    p48_temp1__317 <= p47_temp1__317;
    p48_temp1__318 <= p48_temp1__318_comb;
    p48_temp1__319 <= p47_temp1__319;
    p48_temp1__351 <= p48_temp1__351_comb;
    p48_temp1__344 <= p47_temp1__344;
  end

  // ===== Pipe stage 49:
  wire [31:0] p49_temp1__224_comb;
  wire [31:0] p49_e__56_comb;
  wire [5:0] p49_S1__287_comb;
  wire [4:0] p49_S1__286_comb;
  wire [13:0] p49_S1__285_comb;
  wire [6:0] p49_S1__284_comb;
  wire [1:0] p49_S0__283_comb;
  wire [10:0] p49_S0__282_comb;
  wire [8:0] p49_S0__281_comb;
  wire [9:0] p49_S0__280_comb;
  wire [31:0] p49_and_63299_comb;
  wire [31:0] p49_S1__56_comb;
  wire [31:0] p49_ch__56_comb;
  wire [31:0] p49_S0__55_comb;
  wire [31:0] p49_maj__55_comb;
  wire [31:0] p49_temp1__362_comb;
  wire [31:0] p49_temp1__363_comb;
  wire [31:0] p49_temp2__55_comb;
  wire [31:0] p49_temp1__364_comb;
  wire [31:0] p49_a__56_comb;
  assign p49_temp1__224_comb = p48_temp1__222 + p48_temp1__313;
  assign p49_e__56_comb = p48_a__52 + p49_temp1__224_comb;
  assign p49_S1__287_comb = p49_e__56_comb[5:0] ^ p49_e__56_comb[10:5] ^ p49_e__56_comb[24:19];
  assign p49_S1__286_comb = p49_e__56_comb[31:27] ^ p49_e__56_comb[4:0] ^ p49_e__56_comb[18:14];
  assign p49_S1__285_comb = p49_e__56_comb[26:13] ^ p49_e__56_comb[31:18] ^ p49_e__56_comb[13:0];
  assign p49_S1__284_comb = p49_e__56_comb[12:6] ^ p49_e__56_comb[17:11] ^ p49_e__56_comb[31:25];
  assign p49_S0__283_comb = p48_a__55[1:0] ^ p48_a__55[12:11] ^ p48_a__55[21:20];
  assign p49_S0__282_comb = p48_a__55[31:21] ^ p48_a__55[10:0] ^ p48_a__55[19:9];
  assign p49_S0__281_comb = p48_a__55[20:12] ^ p48_a__55[31:23] ^ p48_a__55[8:0];
  assign p49_S0__280_comb = p48_a__55[11:2] ^ p48_a__55[22:13] ^ p48_a__55[31:22];
  assign p49_and_63299_comb = p48_a__55 & p48_a__54;
  assign p49_S1__56_comb = {p49_S1__287_comb, p49_S1__286_comb, p49_S1__285_comb, p49_S1__284_comb};
  assign p49_ch__56_comb = p49_e__56_comb & p48_e__55 ^ ~(p49_e__56_comb | ~p48_e__54);
  assign p49_S0__55_comb = {p49_S0__283_comb, p49_S0__282_comb, p49_S0__281_comb, p49_S0__280_comb};
  assign p49_maj__55_comb = p49_and_63299_comb ^ p48_a__55 & p48_a__53 ^ p48_and_63174;
  assign p49_temp1__362_comb = p48_e__53 + p49_S1__56_comb;
  assign p49_temp1__363_comb = p49_ch__56_comb + p48_temp1__314;
  assign p49_temp2__55_comb = p49_S0__55_comb + p49_maj__55_comb;
  assign p49_temp1__364_comb = p49_temp1__362_comb + p49_temp1__363_comb;
  assign p49_a__56_comb = p49_temp1__224_comb + p49_temp2__55_comb;

  // Registers for pipe stage 49:
  reg [31:0] p49_value__93;
  reg [31:0] p49_value__96;
  reg [31:0] p49_e__54;
  reg [31:0] p49_e__55;
  reg [31:0] p49_a__53;
  reg [31:0] p49_e__56;
  reg [31:0] p49_a__54;
  reg [31:0] p49_temp1__364;
  reg [31:0] p49_a__55;
  reg [31:0] p49_and_63299;
  reg [31:0] p49_temp1__315;
  reg [31:0] p49_a__56;
  reg [31:0] p49_temp1__316;
  reg [31:0] p49_temp1__317;
  reg [31:0] p49_temp1__318;
  reg [31:0] p49_temp1__319;
  reg [31:0] p49_temp1__351;
  reg [31:0] p49_temp1__344;
  always_ff @ (posedge clk) begin
    p49_value__93 <= p48_value__93;
    p49_value__96 <= p48_value__96;
    p49_e__54 <= p48_e__54;
    p49_e__55 <= p48_e__55;
    p49_a__53 <= p48_a__53;
    p49_e__56 <= p49_e__56_comb;
    p49_a__54 <= p48_a__54;
    p49_temp1__364 <= p49_temp1__364_comb;
    p49_a__55 <= p48_a__55;
    p49_and_63299 <= p49_and_63299_comb;
    p49_temp1__315 <= p48_temp1__315;
    p49_a__56 <= p49_a__56_comb;
    p49_temp1__316 <= p48_temp1__316;
    p49_temp1__317 <= p48_temp1__317;
    p49_temp1__318 <= p48_temp1__318;
    p49_temp1__319 <= p48_temp1__319;
    p49_temp1__351 <= p48_temp1__351;
    p49_temp1__344 <= p48_temp1__344;
  end

  // ===== Pipe stage 50:
  wire [31:0] p50_e__57_comb;
  wire [5:0] p50_S1__291_comb;
  wire [4:0] p50_S1__290_comb;
  wire [13:0] p50_S1__289_comb;
  wire [6:0] p50_S1__288_comb;
  wire [31:0] p50_S1__57_comb;
  wire [1:0] p50_S0__287_comb;
  wire [10:0] p50_S0__286_comb;
  wire [8:0] p50_S0__285_comb;
  wire [9:0] p50_S0__284_comb;
  wire [31:0] p50_and_63382_comb;
  wire [31:0] p50_temp1__229_comb;
  wire [31:0] p50_ch__57_comb;
  wire [31:0] p50_S0__56_comb;
  wire [31:0] p50_maj__56_comb;
  wire [31:0] p50_temp1__230_comb;
  wire [31:0] p50_temp2__56_comb;
  wire [31:0] p50_temp1__232_comb;
  wire [31:0] p50_a__57_comb;
  assign p50_e__57_comb = p49_a__53 + p49_temp1__364;
  assign p50_S1__291_comb = p50_e__57_comb[5:0] ^ p50_e__57_comb[10:5] ^ p50_e__57_comb[24:19];
  assign p50_S1__290_comb = p50_e__57_comb[31:27] ^ p50_e__57_comb[4:0] ^ p50_e__57_comb[18:14];
  assign p50_S1__289_comb = p50_e__57_comb[26:13] ^ p50_e__57_comb[31:18] ^ p50_e__57_comb[13:0];
  assign p50_S1__288_comb = p50_e__57_comb[12:6] ^ p50_e__57_comb[17:11] ^ p50_e__57_comb[31:25];
  assign p50_S1__57_comb = {p50_S1__291_comb, p50_S1__290_comb, p50_S1__289_comb, p50_S1__288_comb};
  assign p50_S0__287_comb = p49_a__56[1:0] ^ p49_a__56[12:11] ^ p49_a__56[21:20];
  assign p50_S0__286_comb = p49_a__56[31:21] ^ p49_a__56[10:0] ^ p49_a__56[19:9];
  assign p50_S0__285_comb = p49_a__56[20:12] ^ p49_a__56[31:23] ^ p49_a__56[8:0];
  assign p50_S0__284_comb = p49_a__56[11:2] ^ p49_a__56[22:13] ^ p49_a__56[31:22];
  assign p50_and_63382_comb = p49_a__56 & p49_a__55;
  assign p50_temp1__229_comb = p49_e__54 + p50_S1__57_comb;
  assign p50_ch__57_comb = p50_e__57_comb & p49_e__56 ^ ~(p50_e__57_comb | ~p49_e__55);
  assign p50_S0__56_comb = {p50_S0__287_comb, p50_S0__286_comb, p50_S0__285_comb, p50_S0__284_comb};
  assign p50_maj__56_comb = p50_and_63382_comb ^ p49_a__56 & p49_a__54 ^ p49_and_63299;
  assign p50_temp1__230_comb = p50_temp1__229_comb + p50_ch__57_comb;
  assign p50_temp2__56_comb = p50_S0__56_comb + p50_maj__56_comb;
  assign p50_temp1__232_comb = p50_temp1__230_comb + p49_temp1__315;
  assign p50_a__57_comb = p49_temp1__364 + p50_temp2__56_comb;

  // Registers for pipe stage 50:
  reg [31:0] p50_value__93;
  reg [31:0] p50_value__96;
  reg [31:0] p50_e__55;
  reg [31:0] p50_e__56;
  reg [31:0] p50_a__54;
  reg [31:0] p50_e__57;
  reg [31:0] p50_a__55;
  reg [31:0] p50_temp1__232;
  reg [31:0] p50_a__56;
  reg [31:0] p50_and_63382;
  reg [31:0] p50_temp1__316;
  reg [31:0] p50_a__57;
  reg [31:0] p50_temp1__317;
  reg [31:0] p50_temp1__318;
  reg [31:0] p50_temp1__319;
  reg [31:0] p50_temp1__351;
  reg [31:0] p50_temp1__344;
  always_ff @ (posedge clk) begin
    p50_value__93 <= p49_value__93;
    p50_value__96 <= p49_value__96;
    p50_e__55 <= p49_e__55;
    p50_e__56 <= p49_e__56;
    p50_a__54 <= p49_a__54;
    p50_e__57 <= p50_e__57_comb;
    p50_a__55 <= p49_a__55;
    p50_temp1__232 <= p50_temp1__232_comb;
    p50_a__56 <= p49_a__56;
    p50_and_63382 <= p50_and_63382_comb;
    p50_temp1__316 <= p49_temp1__316;
    p50_a__57 <= p50_a__57_comb;
    p50_temp1__317 <= p49_temp1__317;
    p50_temp1__318 <= p49_temp1__318;
    p50_temp1__319 <= p49_temp1__319;
    p50_temp1__351 <= p49_temp1__351;
    p50_temp1__344 <= p49_temp1__344;
  end

  // ===== Pipe stage 51:
  wire [1:0] p51_S0__291_comb;
  wire [10:0] p51_S0__290_comb;
  wire [8:0] p51_S0__289_comb;
  wire [9:0] p51_S0__288_comb;
  wire [31:0] p51_and_63464_comb;
  wire [31:0] p51_S0__57_comb;
  wire [31:0] p51_maj__57_comb;
  wire [31:0] p51_e__58_comb;
  wire [31:0] p51_temp2__57_comb;
  wire [31:0] p51_a__58_comb;
  wire [5:0] p51_S1__295_comb;
  wire [4:0] p51_S1__294_comb;
  wire [13:0] p51_S1__293_comb;
  wire [6:0] p51_S1__292_comb;
  wire [31:0] p51_S1__58_comb;
  wire [31:0] p51_ch__58_comb;
  wire [1:0] p51_S0__295_comb;
  wire [10:0] p51_S0__294_comb;
  wire [8:0] p51_S0__293_comb;
  wire [9:0] p51_S0__292_comb;
  wire [31:0] p51_and_63486_comb;
  wire [31:0] p51_temp1__359_comb;
  wire [31:0] p51_temp1__360_comb;
  wire [31:0] p51_S0__58_comb;
  wire [31:0] p51_maj__58_comb;
  wire [31:0] p51_temp1__361_comb;
  wire [31:0] p51_temp2__58_comb;
  wire [31:0] p51_e__59_comb;
  wire [31:0] p51_a__59_comb;
  assign p51_S0__291_comb = p50_a__57[1:0] ^ p50_a__57[12:11] ^ p50_a__57[21:20];
  assign p51_S0__290_comb = p50_a__57[31:21] ^ p50_a__57[10:0] ^ p50_a__57[19:9];
  assign p51_S0__289_comb = p50_a__57[20:12] ^ p50_a__57[31:23] ^ p50_a__57[8:0];
  assign p51_S0__288_comb = p50_a__57[11:2] ^ p50_a__57[22:13] ^ p50_a__57[31:22];
  assign p51_and_63464_comb = p50_a__57 & p50_a__56;
  assign p51_S0__57_comb = {p51_S0__291_comb, p51_S0__290_comb, p51_S0__289_comb, p51_S0__288_comb};
  assign p51_maj__57_comb = p51_and_63464_comb ^ p50_a__57 & p50_a__55 ^ p50_and_63382;
  assign p51_e__58_comb = p50_a__54 + p50_temp1__232;
  assign p51_temp2__57_comb = p51_S0__57_comb + p51_maj__57_comb;
  assign p51_a__58_comb = p50_temp1__232 + p51_temp2__57_comb;
  assign p51_S1__295_comb = p51_e__58_comb[5:0] ^ p51_e__58_comb[10:5] ^ p51_e__58_comb[24:19];
  assign p51_S1__294_comb = p51_e__58_comb[31:27] ^ p51_e__58_comb[4:0] ^ p51_e__58_comb[18:14];
  assign p51_S1__293_comb = p51_e__58_comb[26:13] ^ p51_e__58_comb[31:18] ^ p51_e__58_comb[13:0];
  assign p51_S1__292_comb = p51_e__58_comb[12:6] ^ p51_e__58_comb[17:11] ^ p51_e__58_comb[31:25];
  assign p51_S1__58_comb = {p51_S1__295_comb, p51_S1__294_comb, p51_S1__293_comb, p51_S1__292_comb};
  assign p51_ch__58_comb = p51_e__58_comb & p50_e__57 ^ ~(p51_e__58_comb | ~p50_e__56);
  assign p51_S0__295_comb = p51_a__58_comb[1:0] ^ p51_a__58_comb[12:11] ^ p51_a__58_comb[21:20];
  assign p51_S0__294_comb = p51_a__58_comb[31:21] ^ p51_a__58_comb[10:0] ^ p51_a__58_comb[19:9];
  assign p51_S0__293_comb = p51_a__58_comb[20:12] ^ p51_a__58_comb[31:23] ^ p51_a__58_comb[8:0];
  assign p51_S0__292_comb = p51_a__58_comb[11:2] ^ p51_a__58_comb[22:13] ^ p51_a__58_comb[31:22];
  assign p51_and_63486_comb = p51_a__58_comb & p50_a__57;
  assign p51_temp1__359_comb = p50_e__55 + p51_S1__58_comb;
  assign p51_temp1__360_comb = p51_ch__58_comb + p50_temp1__316;
  assign p51_S0__58_comb = {p51_S0__295_comb, p51_S0__294_comb, p51_S0__293_comb, p51_S0__292_comb};
  assign p51_maj__58_comb = p51_and_63486_comb ^ p51_a__58_comb & p50_a__56 ^ p51_and_63464_comb;
  assign p51_temp1__361_comb = p51_temp1__359_comb + p51_temp1__360_comb;
  assign p51_temp2__58_comb = p51_S0__58_comb + p51_maj__58_comb;
  assign p51_e__59_comb = p50_a__55 + p51_temp1__361_comb;
  assign p51_a__59_comb = p51_temp1__361_comb + p51_temp2__58_comb;

  // Registers for pipe stage 51:
  reg [31:0] p51_value__93;
  reg [31:0] p51_value__96;
  reg [31:0] p51_e__56;
  reg [31:0] p51_e__57;
  reg [31:0] p51_e__58;
  reg [31:0] p51_a__56;
  reg [31:0] p51_a__57;
  reg [31:0] p51_e__59;
  reg [31:0] p51_temp1__317;
  reg [31:0] p51_a__58;
  reg [31:0] p51_and_63486;
  reg [31:0] p51_temp1__318;
  reg [31:0] p51_a__59;
  reg [31:0] p51_temp1__319;
  reg [31:0] p51_temp1__351;
  reg [31:0] p51_temp1__344;
  always_ff @ (posedge clk) begin
    p51_value__93 <= p50_value__93;
    p51_value__96 <= p50_value__96;
    p51_e__56 <= p50_e__56;
    p51_e__57 <= p50_e__57;
    p51_e__58 <= p51_e__58_comb;
    p51_a__56 <= p50_a__56;
    p51_a__57 <= p50_a__57;
    p51_e__59 <= p51_e__59_comb;
    p51_temp1__317 <= p50_temp1__317;
    p51_a__58 <= p51_a__58_comb;
    p51_and_63486 <= p51_and_63486_comb;
    p51_temp1__318 <= p50_temp1__318;
    p51_a__59 <= p51_a__59_comb;
    p51_temp1__319 <= p50_temp1__319;
    p51_temp1__351 <= p50_temp1__351;
    p51_temp1__344 <= p50_temp1__344;
  end

  // ===== Pipe stage 52:
  wire [5:0] p52_S1__299_comb;
  wire [4:0] p52_S1__298_comb;
  wire [13:0] p52_S1__297_comb;
  wire [6:0] p52_S1__296_comb;
  wire [31:0] p52_S1__59_comb;
  wire [31:0] p52_ch__59_comb;
  wire [31:0] p52_temp1__356_comb;
  wire [31:0] p52_temp1__357_comb;
  wire [31:0] p52_temp1__358_comb;
  wire [31:0] p52_e__60_comb;
  wire [1:0] p52_S0__299_comb;
  wire [10:0] p52_S0__298_comb;
  wire [8:0] p52_S0__297_comb;
  wire [9:0] p52_S0__296_comb;
  wire [31:0] p52_and_63588_comb;
  wire [5:0] p52_S1__303_comb;
  wire [4:0] p52_S1__302_comb;
  wire [13:0] p52_S1__301_comb;
  wire [6:0] p52_S1__300_comb;
  wire [31:0] p52_S0__59_comb;
  wire [31:0] p52_maj__59_comb;
  wire [31:0] p52_S1__60_comb;
  wire [31:0] p52_ch__60_comb;
  wire [31:0] p52_temp2__59_comb;
  wire [31:0] p52_temp1__353_comb;
  wire [31:0] p52_temp1__354_comb;
  wire [31:0] p52_a__60_comb;
  assign p52_S1__299_comb = p51_e__59[5:0] ^ p51_e__59[10:5] ^ p51_e__59[24:19];
  assign p52_S1__298_comb = p51_e__59[31:27] ^ p51_e__59[4:0] ^ p51_e__59[18:14];
  assign p52_S1__297_comb = p51_e__59[26:13] ^ p51_e__59[31:18] ^ p51_e__59[13:0];
  assign p52_S1__296_comb = p51_e__59[12:6] ^ p51_e__59[17:11] ^ p51_e__59[31:25];
  assign p52_S1__59_comb = {p52_S1__299_comb, p52_S1__298_comb, p52_S1__297_comb, p52_S1__296_comb};
  assign p52_ch__59_comb = p51_e__59 & p51_e__58 ^ ~(p51_e__59 | ~p51_e__57);
  assign p52_temp1__356_comb = p51_e__56 + p52_S1__59_comb;
  assign p52_temp1__357_comb = p52_ch__59_comb + p51_temp1__317;
  assign p52_temp1__358_comb = p52_temp1__356_comb + p52_temp1__357_comb;
  assign p52_e__60_comb = p51_a__56 + p52_temp1__358_comb;
  assign p52_S0__299_comb = p51_a__59[1:0] ^ p51_a__59[12:11] ^ p51_a__59[21:20];
  assign p52_S0__298_comb = p51_a__59[31:21] ^ p51_a__59[10:0] ^ p51_a__59[19:9];
  assign p52_S0__297_comb = p51_a__59[20:12] ^ p51_a__59[31:23] ^ p51_a__59[8:0];
  assign p52_S0__296_comb = p51_a__59[11:2] ^ p51_a__59[22:13] ^ p51_a__59[31:22];
  assign p52_and_63588_comb = p51_a__59 & p51_a__58;
  assign p52_S1__303_comb = p52_e__60_comb[5:0] ^ p52_e__60_comb[10:5] ^ p52_e__60_comb[24:19];
  assign p52_S1__302_comb = p52_e__60_comb[31:27] ^ p52_e__60_comb[4:0] ^ p52_e__60_comb[18:14];
  assign p52_S1__301_comb = p52_e__60_comb[26:13] ^ p52_e__60_comb[31:18] ^ p52_e__60_comb[13:0];
  assign p52_S1__300_comb = p52_e__60_comb[12:6] ^ p52_e__60_comb[17:11] ^ p52_e__60_comb[31:25];
  assign p52_S0__59_comb = {p52_S0__299_comb, p52_S0__298_comb, p52_S0__297_comb, p52_S0__296_comb};
  assign p52_maj__59_comb = p52_and_63588_comb ^ p51_a__59 & p51_a__57 ^ p51_and_63486;
  assign p52_S1__60_comb = {p52_S1__303_comb, p52_S1__302_comb, p52_S1__301_comb, p52_S1__300_comb};
  assign p52_ch__60_comb = p52_e__60_comb & p51_e__59 ^ ~(p52_e__60_comb | ~p51_e__58);
  assign p52_temp2__59_comb = p52_S0__59_comb + p52_maj__59_comb;
  assign p52_temp1__353_comb = p51_e__57 + p52_S1__60_comb;
  assign p52_temp1__354_comb = p52_ch__60_comb + p51_temp1__318;
  assign p52_a__60_comb = p52_temp1__358_comb + p52_temp2__59_comb;

  // Registers for pipe stage 52:
  reg [31:0] p52_value__93;
  reg [31:0] p52_value__96;
  reg [31:0] p52_e__58;
  reg [31:0] p52_a__57;
  reg [31:0] p52_e__59;
  reg [31:0] p52_a__58;
  reg [31:0] p52_e__60;
  reg [31:0] p52_a__59;
  reg [31:0] p52_temp1__353;
  reg [31:0] p52_temp1__354;
  reg [31:0] p52_and_63588;
  reg [31:0] p52_a__60;
  reg [31:0] p52_temp1__319;
  reg [31:0] p52_temp1__351;
  reg [31:0] p52_temp1__344;
  always_ff @ (posedge clk) begin
    p52_value__93 <= p51_value__93;
    p52_value__96 <= p51_value__96;
    p52_e__58 <= p51_e__58;
    p52_a__57 <= p51_a__57;
    p52_e__59 <= p51_e__59;
    p52_a__58 <= p51_a__58;
    p52_e__60 <= p52_e__60_comb;
    p52_a__59 <= p51_a__59;
    p52_temp1__353 <= p52_temp1__353_comb;
    p52_temp1__354 <= p52_temp1__354_comb;
    p52_and_63588 <= p52_and_63588_comb;
    p52_a__60 <= p52_a__60_comb;
    p52_temp1__319 <= p51_temp1__319;
    p52_temp1__351 <= p51_temp1__351;
    p52_temp1__344 <= p51_temp1__344;
  end

  // ===== Pipe stage 53:
  wire [31:0] p53_temp1__355_comb;
  wire [31:0] p53_e__61_comb;
  wire [5:0] p53_S1__307_comb;
  wire [4:0] p53_S1__306_comb;
  wire [13:0] p53_S1__305_comb;
  wire [6:0] p53_S1__304_comb;
  wire [1:0] p53_S0__303_comb;
  wire [10:0] p53_S0__302_comb;
  wire [8:0] p53_S0__301_comb;
  wire [9:0] p53_S0__300_comb;
  wire [31:0] p53_and_63662_comb;
  wire [31:0] p53_S1__61_comb;
  wire [31:0] p53_S0__60_comb;
  wire [31:0] p53_maj__60_comb;
  wire [31:0] p53_temp1__245_comb;
  wire [31:0] p53_ch__61_comb;
  wire [31:0] p53_temp2__60_comb;
  wire [31:0] p53_temp1__246_comb;
  wire [31:0] p53_a__61_comb;
  assign p53_temp1__355_comb = p52_temp1__353 + p52_temp1__354;
  assign p53_e__61_comb = p52_a__57 + p53_temp1__355_comb;
  assign p53_S1__307_comb = p53_e__61_comb[5:0] ^ p53_e__61_comb[10:5] ^ p53_e__61_comb[24:19];
  assign p53_S1__306_comb = p53_e__61_comb[31:27] ^ p53_e__61_comb[4:0] ^ p53_e__61_comb[18:14];
  assign p53_S1__305_comb = p53_e__61_comb[26:13] ^ p53_e__61_comb[31:18] ^ p53_e__61_comb[13:0];
  assign p53_S1__304_comb = p53_e__61_comb[12:6] ^ p53_e__61_comb[17:11] ^ p53_e__61_comb[31:25];
  assign p53_S0__303_comb = p52_a__60[1:0] ^ p52_a__60[12:11] ^ p52_a__60[21:20];
  assign p53_S0__302_comb = p52_a__60[31:21] ^ p52_a__60[10:0] ^ p52_a__60[19:9];
  assign p53_S0__301_comb = p52_a__60[20:12] ^ p52_a__60[31:23] ^ p52_a__60[8:0];
  assign p53_S0__300_comb = p52_a__60[11:2] ^ p52_a__60[22:13] ^ p52_a__60[31:22];
  assign p53_and_63662_comb = p52_a__60 & p52_a__59;
  assign p53_S1__61_comb = {p53_S1__307_comb, p53_S1__306_comb, p53_S1__305_comb, p53_S1__304_comb};
  assign p53_S0__60_comb = {p53_S0__303_comb, p53_S0__302_comb, p53_S0__301_comb, p53_S0__300_comb};
  assign p53_maj__60_comb = p53_and_63662_comb ^ p52_a__60 & p52_a__58 ^ p52_and_63588;
  assign p53_temp1__245_comb = p52_e__58 + p53_S1__61_comb;
  assign p53_ch__61_comb = p53_e__61_comb & p52_e__60 ^ ~(p53_e__61_comb | ~p52_e__59);
  assign p53_temp2__60_comb = p53_S0__60_comb + p53_maj__60_comb;
  assign p53_temp1__246_comb = p53_temp1__245_comb + p53_ch__61_comb;
  assign p53_a__61_comb = p53_temp1__355_comb + p53_temp2__60_comb;

  // Registers for pipe stage 53:
  reg [31:0] p53_value__93;
  reg [31:0] p53_value__96;
  reg [31:0] p53_e__59;
  reg [31:0] p53_a__58;
  reg [31:0] p53_e__60;
  reg [31:0] p53_a__59;
  reg [31:0] p53_e__61;
  reg [31:0] p53_a__60;
  reg [31:0] p53_and_63662;
  reg [31:0] p53_temp1__246;
  reg [31:0] p53_temp1__319;
  reg [31:0] p53_a__61;
  reg [31:0] p53_temp1__351;
  reg [31:0] p53_temp1__344;
  always_ff @ (posedge clk) begin
    p53_value__93 <= p52_value__93;
    p53_value__96 <= p52_value__96;
    p53_e__59 <= p52_e__59;
    p53_a__58 <= p52_a__58;
    p53_e__60 <= p52_e__60;
    p53_a__59 <= p52_a__59;
    p53_e__61 <= p53_e__61_comb;
    p53_a__60 <= p52_a__60;
    p53_and_63662 <= p53_and_63662_comb;
    p53_temp1__246 <= p53_temp1__246_comb;
    p53_temp1__319 <= p52_temp1__319;
    p53_a__61 <= p53_a__61_comb;
    p53_temp1__351 <= p52_temp1__351;
    p53_temp1__344 <= p52_temp1__344;
  end

  // ===== Pipe stage 54:
  wire [31:0] p54_temp1__248_comb;
  wire [31:0] p54_e__62_comb;
  wire [5:0] p54_S1__311_comb;
  wire [4:0] p54_S1__310_comb;
  wire [13:0] p54_S1__309_comb;
  wire [6:0] p54_S1__308_comb;
  wire [1:0] p54_S0__307_comb;
  wire [10:0] p54_S0__306_comb;
  wire [8:0] p54_S0__305_comb;
  wire [9:0] p54_S0__304_comb;
  wire [31:0] p54_and_63730_comb;
  wire [31:0] p54_S1__62_comb;
  wire [31:0] p54_ch__62_comb;
  wire [31:0] p54_S0__61_comb;
  wire [31:0] p54_maj__61_comb;
  wire [31:0] p54_temp1__346_comb;
  wire [31:0] p54_temp1__347_comb;
  wire [31:0] p54_temp2__61_comb;
  wire [31:0] p54_temp1__350_comb;
  wire [31:0] p54_a__62_comb;
  assign p54_temp1__248_comb = p53_temp1__246 + p53_temp1__319;
  assign p54_e__62_comb = p53_a__58 + p54_temp1__248_comb;
  assign p54_S1__311_comb = p54_e__62_comb[5:0] ^ p54_e__62_comb[10:5] ^ p54_e__62_comb[24:19];
  assign p54_S1__310_comb = p54_e__62_comb[31:27] ^ p54_e__62_comb[4:0] ^ p54_e__62_comb[18:14];
  assign p54_S1__309_comb = p54_e__62_comb[26:13] ^ p54_e__62_comb[31:18] ^ p54_e__62_comb[13:0];
  assign p54_S1__308_comb = p54_e__62_comb[12:6] ^ p54_e__62_comb[17:11] ^ p54_e__62_comb[31:25];
  assign p54_S0__307_comb = p53_a__61[1:0] ^ p53_a__61[12:11] ^ p53_a__61[21:20];
  assign p54_S0__306_comb = p53_a__61[31:21] ^ p53_a__61[10:0] ^ p53_a__61[19:9];
  assign p54_S0__305_comb = p53_a__61[20:12] ^ p53_a__61[31:23] ^ p53_a__61[8:0];
  assign p54_S0__304_comb = p53_a__61[11:2] ^ p53_a__61[22:13] ^ p53_a__61[31:22];
  assign p54_and_63730_comb = p53_a__61 & p53_a__60;
  assign p54_S1__62_comb = {p54_S1__311_comb, p54_S1__310_comb, p54_S1__309_comb, p54_S1__308_comb};
  assign p54_ch__62_comb = p54_e__62_comb & p53_e__61 ^ ~(p54_e__62_comb | ~p53_e__60);
  assign p54_S0__61_comb = {p54_S0__307_comb, p54_S0__306_comb, p54_S0__305_comb, p54_S0__304_comb};
  assign p54_maj__61_comb = p54_and_63730_comb ^ p53_a__61 & p53_a__59 ^ p53_and_63662;
  assign p54_temp1__346_comb = p53_e__59 + p54_S1__62_comb;
  assign p54_temp1__347_comb = p54_ch__62_comb + p53_value__93;
  assign p54_temp2__61_comb = p54_S0__61_comb + p54_maj__61_comb;
  assign p54_temp1__350_comb = p54_temp1__346_comb + p54_temp1__347_comb;
  assign p54_a__62_comb = p54_temp1__248_comb + p54_temp2__61_comb;

  // Registers for pipe stage 54:
  reg [31:0] p54_value__96;
  reg [31:0] p54_e__60;
  reg [31:0] p54_a__59;
  reg [31:0] p54_e__61;
  reg [31:0] p54_a__60;
  reg [31:0] p54_e__62;
  reg [31:0] p54_a__61;
  reg [31:0] p54_and_63730;
  reg [31:0] p54_temp1__350;
  reg [31:0] p54_temp1__351;
  reg [31:0] p54_a__62;
  reg [31:0] p54_temp1__344;
  always_ff @ (posedge clk) begin
    p54_value__96 <= p53_value__96;
    p54_e__60 <= p53_e__60;
    p54_a__59 <= p53_a__59;
    p54_e__61 <= p53_e__61;
    p54_a__60 <= p53_a__60;
    p54_e__62 <= p54_e__62_comb;
    p54_a__61 <= p53_a__61;
    p54_and_63730 <= p54_and_63730_comb;
    p54_temp1__350 <= p54_temp1__350_comb;
    p54_temp1__351 <= p53_temp1__351;
    p54_a__62 <= p54_a__62_comb;
    p54_temp1__344 <= p53_temp1__344;
  end

  // ===== Pipe stage 55:
  wire [31:0] p55_temp1__352_comb;
  wire [1:0] p55_S0__311_comb;
  wire [10:0] p55_S0__310_comb;
  wire [8:0] p55_S0__309_comb;
  wire [9:0] p55_S0__308_comb;
  wire [31:0] p55_and_63788_comb;
  wire [31:0] p55_e__63_comb;
  wire [31:0] p55_S0__62_comb;
  wire [31:0] p55_maj__62_comb;
  wire [31:0] p55_temp2__62_comb;
  wire [5:0] p55_S1__315_comb;
  wire [4:0] p55_S1__314_comb;
  wire [13:0] p55_S1__313_comb;
  wire [6:0] p55_S1__312_comb;
  wire [31:0] p55_a__63_comb;
  wire [31:0] p55_S1__63_comb;
  wire [31:0] p55_ch__63_comb;
  wire [31:0] p55_temp1__339_comb;
  wire [31:0] p55_temp1__340_comb;
  wire [30:0] p55_add_63830_comb;
  wire [30:0] p55_add_63832_comb;
  wire [29:0] p55_add_63834_comb;
  wire [31:0] p55_h__1_comb;
  wire [31:0] p55_h7_comb;
  wire [31:0] p55_maj__63_comb;
  wire [31:0] p55_b__4_comb;
  wire [31:0] p55_temp1__343_comb;
  wire [31:0] p55_concat_63838_comb;
  wire [31:0] p55_concat_63839_comb;
  wire [31:0] p55_concat_63840_comb;
  wire [31:0] p55_add_63841_comb;
  wire [31:0] p55_add_63842_comb;
  wire [31:0] p55_add_63829_comb;
  assign p55_temp1__352_comb = p54_temp1__350 + p54_temp1__351;
  assign p55_S0__311_comb = p54_a__62[1:0] ^ p54_a__62[12:11] ^ p54_a__62[21:20];
  assign p55_S0__310_comb = p54_a__62[31:21] ^ p54_a__62[10:0] ^ p54_a__62[19:9];
  assign p55_S0__309_comb = p54_a__62[20:12] ^ p54_a__62[31:23] ^ p54_a__62[8:0];
  assign p55_S0__308_comb = p54_a__62[11:2] ^ p54_a__62[22:13] ^ p54_a__62[31:22];
  assign p55_and_63788_comb = p54_a__62 & p54_a__61;
  assign p55_e__63_comb = p54_a__59 + p55_temp1__352_comb;
  assign p55_S0__62_comb = {p55_S0__311_comb, p55_S0__310_comb, p55_S0__309_comb, p55_S0__308_comb};
  assign p55_maj__62_comb = p55_and_63788_comb ^ p54_a__62 & p54_a__60 ^ p54_and_63730;
  assign p55_temp2__62_comb = p55_S0__62_comb + p55_maj__62_comb;
  assign p55_S1__315_comb = p55_e__63_comb[5:0] ^ p55_e__63_comb[10:5] ^ p55_e__63_comb[24:19];
  assign p55_S1__314_comb = p55_e__63_comb[31:27] ^ p55_e__63_comb[4:0] ^ p55_e__63_comb[18:14];
  assign p55_S1__313_comb = p55_e__63_comb[26:13] ^ p55_e__63_comb[31:18] ^ p55_e__63_comb[13:0];
  assign p55_S1__312_comb = p55_e__63_comb[12:6] ^ p55_e__63_comb[17:11] ^ p55_e__63_comb[31:25];
  assign p55_a__63_comb = p55_temp1__352_comb + p55_temp2__62_comb;
  assign p55_S1__63_comb = {p55_S1__315_comb, p55_S1__314_comb, p55_S1__313_comb, p55_S1__312_comb};
  assign p55_ch__63_comb = p55_e__63_comb & p54_e__62 ^ ~(p55_e__63_comb | ~p54_e__61);
  assign p55_temp1__339_comb = p54_e__60 + p55_S1__63_comb;
  assign p55_temp1__340_comb = p55_ch__63_comb + p54_value__96;
  assign p55_add_63830_comb = p54_a__62[31:1] + 31'h1e37_79b9;
  assign p55_add_63832_comb = p54_a__61[31:1] + 31'h52a7_fa9d;
  assign p55_add_63834_comb = p55_e__63_comb[31:2] + 30'h26c1_5a23;
  assign p55_h__1_comb = 32'h1f83_d9ab;
  assign p55_h7_comb = 32'h5be0_cd19;
  assign p55_maj__63_comb = p55_a__63_comb & p54_a__62 ^ p55_a__63_comb & p54_a__61 ^ p55_and_63788_comb;
  assign p55_b__4_comb = 32'h6a09_e667;
  assign p55_temp1__343_comb = p55_temp1__339_comb + p55_temp1__340_comb;
  assign p55_concat_63838_comb = {p55_add_63830_comb, p54_a__62[0]};
  assign p55_concat_63839_comb = {p55_add_63832_comb, p54_a__61[0]};
  assign p55_concat_63840_comb = {p55_add_63834_comb, p55_e__63_comb[1:0]};
  assign p55_add_63841_comb = p54_e__62 + p55_h__1_comb;
  assign p55_add_63842_comb = p54_e__61 + p55_h7_comb;
  assign p55_add_63829_comb = p55_maj__63_comb + p55_b__4_comb;

  // Registers for pipe stage 55:
  reg [31:0] p55_a__60;
  reg [31:0] p55_a__63;
  reg [31:0] p55_temp1__343;
  reg [31:0] p55_temp1__344;
  reg [31:0] p55_concat_63838;
  reg [31:0] p55_concat_63839;
  reg [31:0] p55_concat_63840;
  reg [31:0] p55_add_63841;
  reg [31:0] p55_add_63842;
  reg [31:0] p55_add_63829;
  always_ff @ (posedge clk) begin
    p55_a__60 <= p54_a__60;
    p55_a__63 <= p55_a__63_comb;
    p55_temp1__343 <= p55_temp1__343_comb;
    p55_temp1__344 <= p54_temp1__344;
    p55_concat_63838 <= p55_concat_63838_comb;
    p55_concat_63839 <= p55_concat_63839_comb;
    p55_concat_63840 <= p55_concat_63840_comb;
    p55_add_63841 <= p55_add_63841_comb;
    p55_add_63842 <= p55_add_63842_comb;
    p55_add_63829 <= p55_add_63829_comb;
  end

  // ===== Pipe stage 56:
  wire [1:0] p56_S0__315_comb;
  wire [10:0] p56_S0__314_comb;
  wire [8:0] p56_S0__313_comb;
  wire [9:0] p56_S0__312_comb;
  wire [31:0] p56_S0__63_comb;
  wire [31:0] p56_temp1__345_comb;
  wire [31:0] p56_add_63881_comb;
  wire [31:0] p56_c__2_comb;
  wire [31:0] p56_e__64_comb;
  wire [31:0] p56_f__2_comb;
  wire [31:0] p56_add_63885_comb;
  wire [31:0] p56_add_63886_comb;
  wire [31:0] p56_add_63887_comb;
  wire [255:0] p56_tuple_63888_comb;
  assign p56_S0__315_comb = p55_a__63[1:0] ^ p55_a__63[12:11] ^ p55_a__63[21:20];
  assign p56_S0__314_comb = p55_a__63[31:21] ^ p55_a__63[10:0] ^ p55_a__63[19:9];
  assign p56_S0__313_comb = p55_a__63[20:12] ^ p55_a__63[31:23] ^ p55_a__63[8:0];
  assign p56_S0__312_comb = p55_a__63[11:2] ^ p55_a__63[22:13] ^ p55_a__63[31:22];
  assign p56_S0__63_comb = {p56_S0__315_comb, p56_S0__314_comb, p56_S0__313_comb, p56_S0__312_comb};
  assign p56_temp1__345_comb = p55_temp1__343 + p55_temp1__344;
  assign p56_add_63881_comb = p56_S0__63_comb + p56_temp1__345_comb;
  assign p56_c__2_comb = 32'hbb67_ae85;
  assign p56_e__64_comb = p55_a__60 + p56_temp1__345_comb;
  assign p56_f__2_comb = 32'h510e_527f;
  assign p56_add_63885_comb = p56_add_63881_comb + p55_add_63829;
  assign p56_add_63886_comb = p55_a__63 + p56_c__2_comb;
  assign p56_add_63887_comb = p56_e__64_comb + p56_f__2_comb;
  assign p56_tuple_63888_comb = {p56_add_63885_comb, p56_add_63886_comb, p55_concat_63838, p55_concat_63839, p56_add_63887_comb, p55_concat_63840, p55_add_63841, p55_add_63842};

  // Registers for pipe stage 56:
  reg [255:0] p56_tuple_63888;
  always_ff @ (posedge clk) begin
    p56_tuple_63888 <= p56_tuple_63888_comb;
  end
  assign out = p56_tuple_63888;
endmodule
