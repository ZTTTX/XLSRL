module xls_test(
  input wire clk,
  input wire [2047:0] a,
  input wire [2047:0] b,
  input wire [2047:0] result,
  output wire [6143:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] smul32b_32b_x_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    reg signed [31:0] signed_lhs;
    reg signed [31:0] signed_rhs;
    reg signed [31:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul32b_32b_x_32b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  wire [31:0] a_unflattened[8][8];
  assign a_unflattened[0][0] = a[31:0];
  assign a_unflattened[0][1] = a[63:32];
  assign a_unflattened[0][2] = a[95:64];
  assign a_unflattened[0][3] = a[127:96];
  assign a_unflattened[0][4] = a[159:128];
  assign a_unflattened[0][5] = a[191:160];
  assign a_unflattened[0][6] = a[223:192];
  assign a_unflattened[0][7] = a[255:224];
  assign a_unflattened[1][0] = a[287:256];
  assign a_unflattened[1][1] = a[319:288];
  assign a_unflattened[1][2] = a[351:320];
  assign a_unflattened[1][3] = a[383:352];
  assign a_unflattened[1][4] = a[415:384];
  assign a_unflattened[1][5] = a[447:416];
  assign a_unflattened[1][6] = a[479:448];
  assign a_unflattened[1][7] = a[511:480];
  assign a_unflattened[2][0] = a[543:512];
  assign a_unflattened[2][1] = a[575:544];
  assign a_unflattened[2][2] = a[607:576];
  assign a_unflattened[2][3] = a[639:608];
  assign a_unflattened[2][4] = a[671:640];
  assign a_unflattened[2][5] = a[703:672];
  assign a_unflattened[2][6] = a[735:704];
  assign a_unflattened[2][7] = a[767:736];
  assign a_unflattened[3][0] = a[799:768];
  assign a_unflattened[3][1] = a[831:800];
  assign a_unflattened[3][2] = a[863:832];
  assign a_unflattened[3][3] = a[895:864];
  assign a_unflattened[3][4] = a[927:896];
  assign a_unflattened[3][5] = a[959:928];
  assign a_unflattened[3][6] = a[991:960];
  assign a_unflattened[3][7] = a[1023:992];
  assign a_unflattened[4][0] = a[1055:1024];
  assign a_unflattened[4][1] = a[1087:1056];
  assign a_unflattened[4][2] = a[1119:1088];
  assign a_unflattened[4][3] = a[1151:1120];
  assign a_unflattened[4][4] = a[1183:1152];
  assign a_unflattened[4][5] = a[1215:1184];
  assign a_unflattened[4][6] = a[1247:1216];
  assign a_unflattened[4][7] = a[1279:1248];
  assign a_unflattened[5][0] = a[1311:1280];
  assign a_unflattened[5][1] = a[1343:1312];
  assign a_unflattened[5][2] = a[1375:1344];
  assign a_unflattened[5][3] = a[1407:1376];
  assign a_unflattened[5][4] = a[1439:1408];
  assign a_unflattened[5][5] = a[1471:1440];
  assign a_unflattened[5][6] = a[1503:1472];
  assign a_unflattened[5][7] = a[1535:1504];
  assign a_unflattened[6][0] = a[1567:1536];
  assign a_unflattened[6][1] = a[1599:1568];
  assign a_unflattened[6][2] = a[1631:1600];
  assign a_unflattened[6][3] = a[1663:1632];
  assign a_unflattened[6][4] = a[1695:1664];
  assign a_unflattened[6][5] = a[1727:1696];
  assign a_unflattened[6][6] = a[1759:1728];
  assign a_unflattened[6][7] = a[1791:1760];
  assign a_unflattened[7][0] = a[1823:1792];
  assign a_unflattened[7][1] = a[1855:1824];
  assign a_unflattened[7][2] = a[1887:1856];
  assign a_unflattened[7][3] = a[1919:1888];
  assign a_unflattened[7][4] = a[1951:1920];
  assign a_unflattened[7][5] = a[1983:1952];
  assign a_unflattened[7][6] = a[2015:1984];
  assign a_unflattened[7][7] = a[2047:2016];
  wire [31:0] b_unflattened[8][8];
  assign b_unflattened[0][0] = b[31:0];
  assign b_unflattened[0][1] = b[63:32];
  assign b_unflattened[0][2] = b[95:64];
  assign b_unflattened[0][3] = b[127:96];
  assign b_unflattened[0][4] = b[159:128];
  assign b_unflattened[0][5] = b[191:160];
  assign b_unflattened[0][6] = b[223:192];
  assign b_unflattened[0][7] = b[255:224];
  assign b_unflattened[1][0] = b[287:256];
  assign b_unflattened[1][1] = b[319:288];
  assign b_unflattened[1][2] = b[351:320];
  assign b_unflattened[1][3] = b[383:352];
  assign b_unflattened[1][4] = b[415:384];
  assign b_unflattened[1][5] = b[447:416];
  assign b_unflattened[1][6] = b[479:448];
  assign b_unflattened[1][7] = b[511:480];
  assign b_unflattened[2][0] = b[543:512];
  assign b_unflattened[2][1] = b[575:544];
  assign b_unflattened[2][2] = b[607:576];
  assign b_unflattened[2][3] = b[639:608];
  assign b_unflattened[2][4] = b[671:640];
  assign b_unflattened[2][5] = b[703:672];
  assign b_unflattened[2][6] = b[735:704];
  assign b_unflattened[2][7] = b[767:736];
  assign b_unflattened[3][0] = b[799:768];
  assign b_unflattened[3][1] = b[831:800];
  assign b_unflattened[3][2] = b[863:832];
  assign b_unflattened[3][3] = b[895:864];
  assign b_unflattened[3][4] = b[927:896];
  assign b_unflattened[3][5] = b[959:928];
  assign b_unflattened[3][6] = b[991:960];
  assign b_unflattened[3][7] = b[1023:992];
  assign b_unflattened[4][0] = b[1055:1024];
  assign b_unflattened[4][1] = b[1087:1056];
  assign b_unflattened[4][2] = b[1119:1088];
  assign b_unflattened[4][3] = b[1151:1120];
  assign b_unflattened[4][4] = b[1183:1152];
  assign b_unflattened[4][5] = b[1215:1184];
  assign b_unflattened[4][6] = b[1247:1216];
  assign b_unflattened[4][7] = b[1279:1248];
  assign b_unflattened[5][0] = b[1311:1280];
  assign b_unflattened[5][1] = b[1343:1312];
  assign b_unflattened[5][2] = b[1375:1344];
  assign b_unflattened[5][3] = b[1407:1376];
  assign b_unflattened[5][4] = b[1439:1408];
  assign b_unflattened[5][5] = b[1471:1440];
  assign b_unflattened[5][6] = b[1503:1472];
  assign b_unflattened[5][7] = b[1535:1504];
  assign b_unflattened[6][0] = b[1567:1536];
  assign b_unflattened[6][1] = b[1599:1568];
  assign b_unflattened[6][2] = b[1631:1600];
  assign b_unflattened[6][3] = b[1663:1632];
  assign b_unflattened[6][4] = b[1695:1664];
  assign b_unflattened[6][5] = b[1727:1696];
  assign b_unflattened[6][6] = b[1759:1728];
  assign b_unflattened[6][7] = b[1791:1760];
  assign b_unflattened[7][0] = b[1823:1792];
  assign b_unflattened[7][1] = b[1855:1824];
  assign b_unflattened[7][2] = b[1887:1856];
  assign b_unflattened[7][3] = b[1919:1888];
  assign b_unflattened[7][4] = b[1951:1920];
  assign b_unflattened[7][5] = b[1983:1952];
  assign b_unflattened[7][6] = b[2015:1984];
  assign b_unflattened[7][7] = b[2047:2016];
  wire [31:0] result_unflattened[8][8];
  assign result_unflattened[0][0] = result[31:0];
  assign result_unflattened[0][1] = result[63:32];
  assign result_unflattened[0][2] = result[95:64];
  assign result_unflattened[0][3] = result[127:96];
  assign result_unflattened[0][4] = result[159:128];
  assign result_unflattened[0][5] = result[191:160];
  assign result_unflattened[0][6] = result[223:192];
  assign result_unflattened[0][7] = result[255:224];
  assign result_unflattened[1][0] = result[287:256];
  assign result_unflattened[1][1] = result[319:288];
  assign result_unflattened[1][2] = result[351:320];
  assign result_unflattened[1][3] = result[383:352];
  assign result_unflattened[1][4] = result[415:384];
  assign result_unflattened[1][5] = result[447:416];
  assign result_unflattened[1][6] = result[479:448];
  assign result_unflattened[1][7] = result[511:480];
  assign result_unflattened[2][0] = result[543:512];
  assign result_unflattened[2][1] = result[575:544];
  assign result_unflattened[2][2] = result[607:576];
  assign result_unflattened[2][3] = result[639:608];
  assign result_unflattened[2][4] = result[671:640];
  assign result_unflattened[2][5] = result[703:672];
  assign result_unflattened[2][6] = result[735:704];
  assign result_unflattened[2][7] = result[767:736];
  assign result_unflattened[3][0] = result[799:768];
  assign result_unflattened[3][1] = result[831:800];
  assign result_unflattened[3][2] = result[863:832];
  assign result_unflattened[3][3] = result[895:864];
  assign result_unflattened[3][4] = result[927:896];
  assign result_unflattened[3][5] = result[959:928];
  assign result_unflattened[3][6] = result[991:960];
  assign result_unflattened[3][7] = result[1023:992];
  assign result_unflattened[4][0] = result[1055:1024];
  assign result_unflattened[4][1] = result[1087:1056];
  assign result_unflattened[4][2] = result[1119:1088];
  assign result_unflattened[4][3] = result[1151:1120];
  assign result_unflattened[4][4] = result[1183:1152];
  assign result_unflattened[4][5] = result[1215:1184];
  assign result_unflattened[4][6] = result[1247:1216];
  assign result_unflattened[4][7] = result[1279:1248];
  assign result_unflattened[5][0] = result[1311:1280];
  assign result_unflattened[5][1] = result[1343:1312];
  assign result_unflattened[5][2] = result[1375:1344];
  assign result_unflattened[5][3] = result[1407:1376];
  assign result_unflattened[5][4] = result[1439:1408];
  assign result_unflattened[5][5] = result[1471:1440];
  assign result_unflattened[5][6] = result[1503:1472];
  assign result_unflattened[5][7] = result[1535:1504];
  assign result_unflattened[6][0] = result[1567:1536];
  assign result_unflattened[6][1] = result[1599:1568];
  assign result_unflattened[6][2] = result[1631:1600];
  assign result_unflattened[6][3] = result[1663:1632];
  assign result_unflattened[6][4] = result[1695:1664];
  assign result_unflattened[6][5] = result[1727:1696];
  assign result_unflattened[6][6] = result[1759:1728];
  assign result_unflattened[6][7] = result[1791:1760];
  assign result_unflattened[7][0] = result[1823:1792];
  assign result_unflattened[7][1] = result[1855:1824];
  assign result_unflattened[7][2] = result[1887:1856];
  assign result_unflattened[7][3] = result[1919:1888];
  assign result_unflattened[7][4] = result[1951:1920];
  assign result_unflattened[7][5] = result[1983:1952];
  assign result_unflattened[7][6] = result[2015:1984];
  assign result_unflattened[7][7] = result[2047:2016];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_a[8][8];
  reg [31:0] p0_b[8][8];
  always_ff @ (posedge clk) begin
    p0_a <= a_unflattened;
    p0_b <= b_unflattened;
  end

  // ===== Pipe stage 1:
  wire [31:0] p1_array_index_58980_comb;
  wire [31:0] p1_array_index_58981_comb;
  wire [31:0] p1_array_index_58982_comb;
  wire [31:0] p1_array_index_58983_comb;
  wire [31:0] p1_array_index_58986_comb;
  wire [31:0] p1_array_index_58987_comb;
  wire [31:0] p1_array_index_58988_comb;
  wire [31:0] p1_array_index_58989_comb;
  wire [31:0] p1_array_index_58993_comb;
  wire [31:0] p1_array_index_58994_comb;
  wire [31:0] p1_array_index_58996_comb;
  wire [31:0] p1_array_index_58997_comb;
  wire [31:0] p1_array_index_59001_comb;
  wire [31:0] p1_array_index_59002_comb;
  wire [31:0] p1_array_index_59004_comb;
  wire [31:0] p1_array_index_59005_comb;
  wire [31:0] p1_array_index_59009_comb;
  wire [31:0] p1_array_index_59010_comb;
  wire [31:0] p1_array_index_59012_comb;
  wire [31:0] p1_array_index_59013_comb;
  wire [31:0] p1_array_index_59017_comb;
  wire [31:0] p1_array_index_59018_comb;
  wire [31:0] p1_array_index_59020_comb;
  wire [31:0] p1_array_index_59021_comb;
  wire [31:0] p1_array_index_59025_comb;
  wire [31:0] p1_array_index_59026_comb;
  wire [31:0] p1_array_index_59028_comb;
  wire [31:0] p1_array_index_59029_comb;
  wire [31:0] p1_array_index_59033_comb;
  wire [31:0] p1_array_index_59034_comb;
  wire [31:0] p1_array_index_59036_comb;
  wire [31:0] p1_array_index_59037_comb;
  wire [31:0] p1_array_index_59041_comb;
  wire [31:0] p1_array_index_59042_comb;
  wire [31:0] p1_array_index_59044_comb;
  wire [31:0] p1_array_index_59045_comb;
  wire [31:0] p1_array_index_59049_comb;
  wire [31:0] p1_array_index_59050_comb;
  wire [31:0] p1_array_index_59052_comb;
  wire [31:0] p1_array_index_59053_comb;
  wire [31:0] p1_array_index_59057_comb;
  wire [31:0] p1_array_index_59058_comb;
  wire [31:0] p1_array_index_59060_comb;
  wire [31:0] p1_array_index_59061_comb;
  wire [31:0] p1_array_index_59065_comb;
  wire [31:0] p1_array_index_59066_comb;
  wire [31:0] p1_array_index_59068_comb;
  wire [31:0] p1_array_index_59069_comb;
  wire [31:0] p1_array_index_59073_comb;
  wire [31:0] p1_array_index_59074_comb;
  wire [31:0] p1_array_index_59076_comb;
  wire [31:0] p1_array_index_59077_comb;
  wire [31:0] p1_array_index_59081_comb;
  wire [31:0] p1_array_index_59082_comb;
  wire [31:0] p1_array_index_59084_comb;
  wire [31:0] p1_array_index_59085_comb;
  wire [31:0] p1_array_index_59089_comb;
  wire [31:0] p1_array_index_59090_comb;
  wire [31:0] p1_array_index_59092_comb;
  wire [31:0] p1_array_index_59093_comb;
  wire [31:0] p1_array_index_59097_comb;
  wire [31:0] p1_array_index_59098_comb;
  wire [31:0] p1_array_index_59100_comb;
  wire [31:0] p1_array_index_59101_comb;
  wire [31:0] p1_array_index_58978_comb;
  wire [31:0] p1_array_index_58979_comb;
  wire [31:0] p1_array_index_58984_comb;
  wire [31:0] p1_array_index_58985_comb;
  wire [31:0] p1_array_index_58992_comb;
  wire [31:0] p1_array_index_58995_comb;
  wire [31:0] p1_array_index_59000_comb;
  wire [31:0] p1_array_index_59003_comb;
  wire [31:0] p1_array_index_59008_comb;
  wire [31:0] p1_array_index_59011_comb;
  wire [31:0] p1_array_index_59016_comb;
  wire [31:0] p1_array_index_59019_comb;
  wire [31:0] p1_array_index_59024_comb;
  wire [31:0] p1_array_index_59027_comb;
  wire [31:0] p1_array_index_59032_comb;
  wire [31:0] p1_array_index_59035_comb;
  wire [31:0] p1_array_index_59040_comb;
  wire [31:0] p1_array_index_59043_comb;
  wire [31:0] p1_array_index_59048_comb;
  wire [31:0] p1_array_index_59051_comb;
  wire [31:0] p1_array_index_59056_comb;
  wire [31:0] p1_array_index_59059_comb;
  wire [31:0] p1_array_index_59064_comb;
  wire [31:0] p1_array_index_59067_comb;
  wire [31:0] p1_array_index_59072_comb;
  wire [31:0] p1_array_index_59075_comb;
  wire [31:0] p1_array_index_59080_comb;
  wire [31:0] p1_array_index_59083_comb;
  wire [31:0] p1_array_index_59088_comb;
  wire [31:0] p1_array_index_59091_comb;
  wire [31:0] p1_array_index_59096_comb;
  wire [31:0] p1_array_index_59099_comb;
  wire [31:0] p1_array_index_58976_comb;
  wire [31:0] p1_array_index_58977_comb;
  wire [31:0] p1_array_index_58991_comb;
  wire [31:0] p1_array_index_58999_comb;
  wire [31:0] p1_array_index_59007_comb;
  wire [31:0] p1_array_index_59015_comb;
  wire [31:0] p1_array_index_59023_comb;
  wire [31:0] p1_array_index_59031_comb;
  wire [31:0] p1_array_index_59039_comb;
  wire [31:0] p1_array_index_59047_comb;
  wire [31:0] p1_array_index_59055_comb;
  wire [31:0] p1_array_index_59063_comb;
  wire [31:0] p1_array_index_59071_comb;
  wire [31:0] p1_array_index_59079_comb;
  wire [31:0] p1_array_index_59087_comb;
  wire [31:0] p1_array_index_59095_comb;
  wire [31:0] p1_array_index_58974_comb;
  wire [31:0] p1_array_index_58975_comb;
  wire [31:0] p1_array_index_58990_comb;
  wire [31:0] p1_array_index_58998_comb;
  wire [31:0] p1_array_index_59006_comb;
  wire [31:0] p1_array_index_59014_comb;
  wire [31:0] p1_array_index_59022_comb;
  wire [31:0] p1_array_index_59030_comb;
  wire [31:0] p1_array_index_59038_comb;
  wire [31:0] p1_array_index_59046_comb;
  wire [31:0] p1_array_index_59054_comb;
  wire [31:0] p1_array_index_59062_comb;
  wire [31:0] p1_array_index_59070_comb;
  wire [31:0] p1_array_index_59078_comb;
  wire [31:0] p1_array_index_59086_comb;
  wire [31:0] p1_array_index_59094_comb;
  assign p1_array_index_58980_comb = p0_a[3'h0][3'h2];
  assign p1_array_index_58981_comb = p0_b[3'h2][3'h0];
  assign p1_array_index_58982_comb = p0_a[3'h0][3'h4];
  assign p1_array_index_58983_comb = p0_b[3'h4][3'h0];
  assign p1_array_index_58986_comb = p0_a[3'h0][3'h6];
  assign p1_array_index_58987_comb = p0_b[3'h6][3'h0];
  assign p1_array_index_58988_comb = p0_a[3'h0][3'h7];
  assign p1_array_index_58989_comb = p0_b[3'h7][3'h0];
  assign p1_array_index_58993_comb = p0_b[3'h2][3'h1];
  assign p1_array_index_58994_comb = p0_b[3'h4][3'h1];
  assign p1_array_index_58996_comb = p0_b[3'h6][3'h1];
  assign p1_array_index_58997_comb = p0_b[3'h7][3'h1];
  assign p1_array_index_59001_comb = p0_b[3'h2][3'h2];
  assign p1_array_index_59002_comb = p0_b[3'h4][3'h2];
  assign p1_array_index_59004_comb = p0_b[3'h6][3'h2];
  assign p1_array_index_59005_comb = p0_b[3'h7][3'h2];
  assign p1_array_index_59009_comb = p0_b[3'h2][3'h3];
  assign p1_array_index_59010_comb = p0_b[3'h4][3'h3];
  assign p1_array_index_59012_comb = p0_b[3'h6][3'h3];
  assign p1_array_index_59013_comb = p0_b[3'h7][3'h3];
  assign p1_array_index_59017_comb = p0_b[3'h2][3'h4];
  assign p1_array_index_59018_comb = p0_b[3'h4][3'h4];
  assign p1_array_index_59020_comb = p0_b[3'h6][3'h4];
  assign p1_array_index_59021_comb = p0_b[3'h7][3'h4];
  assign p1_array_index_59025_comb = p0_b[3'h2][3'h5];
  assign p1_array_index_59026_comb = p0_b[3'h4][3'h5];
  assign p1_array_index_59028_comb = p0_b[3'h6][3'h5];
  assign p1_array_index_59029_comb = p0_b[3'h7][3'h5];
  assign p1_array_index_59033_comb = p0_b[3'h2][3'h6];
  assign p1_array_index_59034_comb = p0_b[3'h4][3'h6];
  assign p1_array_index_59036_comb = p0_b[3'h6][3'h6];
  assign p1_array_index_59037_comb = p0_b[3'h7][3'h6];
  assign p1_array_index_59041_comb = p0_b[3'h2][3'h7];
  assign p1_array_index_59042_comb = p0_b[3'h4][3'h7];
  assign p1_array_index_59044_comb = p0_b[3'h6][3'h7];
  assign p1_array_index_59045_comb = p0_b[3'h7][3'h7];
  assign p1_array_index_59049_comb = p0_a[3'h1][3'h2];
  assign p1_array_index_59050_comb = p0_a[3'h1][3'h4];
  assign p1_array_index_59052_comb = p0_a[3'h1][3'h6];
  assign p1_array_index_59053_comb = p0_a[3'h1][3'h7];
  assign p1_array_index_59057_comb = p0_a[3'h2][3'h2];
  assign p1_array_index_59058_comb = p0_a[3'h2][3'h4];
  assign p1_array_index_59060_comb = p0_a[3'h2][3'h6];
  assign p1_array_index_59061_comb = p0_a[3'h2][3'h7];
  assign p1_array_index_59065_comb = p0_a[3'h3][3'h2];
  assign p1_array_index_59066_comb = p0_a[3'h3][3'h4];
  assign p1_array_index_59068_comb = p0_a[3'h3][3'h6];
  assign p1_array_index_59069_comb = p0_a[3'h3][3'h7];
  assign p1_array_index_59073_comb = p0_a[3'h4][3'h2];
  assign p1_array_index_59074_comb = p0_a[3'h4][3'h4];
  assign p1_array_index_59076_comb = p0_a[3'h4][3'h6];
  assign p1_array_index_59077_comb = p0_a[3'h4][3'h7];
  assign p1_array_index_59081_comb = p0_a[3'h5][3'h2];
  assign p1_array_index_59082_comb = p0_a[3'h5][3'h4];
  assign p1_array_index_59084_comb = p0_a[3'h5][3'h6];
  assign p1_array_index_59085_comb = p0_a[3'h5][3'h7];
  assign p1_array_index_59089_comb = p0_a[3'h6][3'h2];
  assign p1_array_index_59090_comb = p0_a[3'h6][3'h4];
  assign p1_array_index_59092_comb = p0_a[3'h6][3'h6];
  assign p1_array_index_59093_comb = p0_a[3'h6][3'h7];
  assign p1_array_index_59097_comb = p0_a[3'h7][3'h2];
  assign p1_array_index_59098_comb = p0_a[3'h7][3'h4];
  assign p1_array_index_59100_comb = p0_a[3'h7][3'h6];
  assign p1_array_index_59101_comb = p0_a[3'h7][3'h7];
  assign p1_array_index_58978_comb = p0_a[3'h0][3'h5];
  assign p1_array_index_58979_comb = p0_b[3'h5][3'h0];
  assign p1_array_index_58984_comb = p0_a[3'h0][3'h3];
  assign p1_array_index_58985_comb = p0_b[3'h3][3'h0];
  assign p1_array_index_58992_comb = p0_b[3'h5][3'h1];
  assign p1_array_index_58995_comb = p0_b[3'h3][3'h1];
  assign p1_array_index_59000_comb = p0_b[3'h5][3'h2];
  assign p1_array_index_59003_comb = p0_b[3'h3][3'h2];
  assign p1_array_index_59008_comb = p0_b[3'h5][3'h3];
  assign p1_array_index_59011_comb = p0_b[3'h3][3'h3];
  assign p1_array_index_59016_comb = p0_b[3'h5][3'h4];
  assign p1_array_index_59019_comb = p0_b[3'h3][3'h4];
  assign p1_array_index_59024_comb = p0_b[3'h5][3'h5];
  assign p1_array_index_59027_comb = p0_b[3'h3][3'h5];
  assign p1_array_index_59032_comb = p0_b[3'h5][3'h6];
  assign p1_array_index_59035_comb = p0_b[3'h3][3'h6];
  assign p1_array_index_59040_comb = p0_b[3'h5][3'h7];
  assign p1_array_index_59043_comb = p0_b[3'h3][3'h7];
  assign p1_array_index_59048_comb = p0_a[3'h1][3'h5];
  assign p1_array_index_59051_comb = p0_a[3'h1][3'h3];
  assign p1_array_index_59056_comb = p0_a[3'h2][3'h5];
  assign p1_array_index_59059_comb = p0_a[3'h2][3'h3];
  assign p1_array_index_59064_comb = p0_a[3'h3][3'h5];
  assign p1_array_index_59067_comb = p0_a[3'h3][3'h3];
  assign p1_array_index_59072_comb = p0_a[3'h4][3'h5];
  assign p1_array_index_59075_comb = p0_a[3'h4][3'h3];
  assign p1_array_index_59080_comb = p0_a[3'h5][3'h5];
  assign p1_array_index_59083_comb = p0_a[3'h5][3'h3];
  assign p1_array_index_59088_comb = p0_a[3'h6][3'h5];
  assign p1_array_index_59091_comb = p0_a[3'h6][3'h3];
  assign p1_array_index_59096_comb = p0_a[3'h7][3'h5];
  assign p1_array_index_59099_comb = p0_a[3'h7][3'h3];
  assign p1_array_index_58976_comb = p0_a[3'h0][3'h0];
  assign p1_array_index_58977_comb = p0_b[3'h0][3'h0];
  assign p1_array_index_58991_comb = p0_b[3'h0][3'h1];
  assign p1_array_index_58999_comb = p0_b[3'h0][3'h2];
  assign p1_array_index_59007_comb = p0_b[3'h0][3'h3];
  assign p1_array_index_59015_comb = p0_b[3'h0][3'h4];
  assign p1_array_index_59023_comb = p0_b[3'h0][3'h5];
  assign p1_array_index_59031_comb = p0_b[3'h0][3'h6];
  assign p1_array_index_59039_comb = p0_b[3'h0][3'h7];
  assign p1_array_index_59047_comb = p0_a[3'h1][3'h0];
  assign p1_array_index_59055_comb = p0_a[3'h2][3'h0];
  assign p1_array_index_59063_comb = p0_a[3'h3][3'h0];
  assign p1_array_index_59071_comb = p0_a[3'h4][3'h0];
  assign p1_array_index_59079_comb = p0_a[3'h5][3'h0];
  assign p1_array_index_59087_comb = p0_a[3'h6][3'h0];
  assign p1_array_index_59095_comb = p0_a[3'h7][3'h0];
  assign p1_array_index_58974_comb = p0_a[3'h0][3'h1];
  assign p1_array_index_58975_comb = p0_b[3'h1][3'h0];
  assign p1_array_index_58990_comb = p0_b[3'h1][3'h1];
  assign p1_array_index_58998_comb = p0_b[3'h1][3'h2];
  assign p1_array_index_59006_comb = p0_b[3'h1][3'h3];
  assign p1_array_index_59014_comb = p0_b[3'h1][3'h4];
  assign p1_array_index_59022_comb = p0_b[3'h1][3'h5];
  assign p1_array_index_59030_comb = p0_b[3'h1][3'h6];
  assign p1_array_index_59038_comb = p0_b[3'h1][3'h7];
  assign p1_array_index_59046_comb = p0_a[3'h1][3'h1];
  assign p1_array_index_59054_comb = p0_a[3'h2][3'h1];
  assign p1_array_index_59062_comb = p0_a[3'h3][3'h1];
  assign p1_array_index_59070_comb = p0_a[3'h4][3'h1];
  assign p1_array_index_59078_comb = p0_a[3'h5][3'h1];
  assign p1_array_index_59086_comb = p0_a[3'h6][3'h1];
  assign p1_array_index_59094_comb = p0_a[3'h7][3'h1];

  // Registers for pipe stage 1:
  reg [31:0] p1_a[8][8];
  reg [31:0] p1_b[8][8];
  reg [31:0] p1_array_index_58980;
  reg [31:0] p1_array_index_58981;
  reg [31:0] p1_array_index_58982;
  reg [31:0] p1_array_index_58983;
  reg [31:0] p1_array_index_58986;
  reg [31:0] p1_array_index_58987;
  reg [31:0] p1_array_index_58988;
  reg [31:0] p1_array_index_58989;
  reg [31:0] p1_array_index_58993;
  reg [31:0] p1_array_index_58994;
  reg [31:0] p1_array_index_58996;
  reg [31:0] p1_array_index_58997;
  reg [31:0] p1_array_index_59001;
  reg [31:0] p1_array_index_59002;
  reg [31:0] p1_array_index_59004;
  reg [31:0] p1_array_index_59005;
  reg [31:0] p1_array_index_59009;
  reg [31:0] p1_array_index_59010;
  reg [31:0] p1_array_index_59012;
  reg [31:0] p1_array_index_59013;
  reg [31:0] p1_array_index_59017;
  reg [31:0] p1_array_index_59018;
  reg [31:0] p1_array_index_59020;
  reg [31:0] p1_array_index_59021;
  reg [31:0] p1_array_index_59025;
  reg [31:0] p1_array_index_59026;
  reg [31:0] p1_array_index_59028;
  reg [31:0] p1_array_index_59029;
  reg [31:0] p1_array_index_59033;
  reg [31:0] p1_array_index_59034;
  reg [31:0] p1_array_index_59036;
  reg [31:0] p1_array_index_59037;
  reg [31:0] p1_array_index_59041;
  reg [31:0] p1_array_index_59042;
  reg [31:0] p1_array_index_59044;
  reg [31:0] p1_array_index_59045;
  reg [31:0] p1_array_index_59049;
  reg [31:0] p1_array_index_59050;
  reg [31:0] p1_array_index_59052;
  reg [31:0] p1_array_index_59053;
  reg [31:0] p1_array_index_59057;
  reg [31:0] p1_array_index_59058;
  reg [31:0] p1_array_index_59060;
  reg [31:0] p1_array_index_59061;
  reg [31:0] p1_array_index_59065;
  reg [31:0] p1_array_index_59066;
  reg [31:0] p1_array_index_59068;
  reg [31:0] p1_array_index_59069;
  reg [31:0] p1_array_index_59073;
  reg [31:0] p1_array_index_59074;
  reg [31:0] p1_array_index_59076;
  reg [31:0] p1_array_index_59077;
  reg [31:0] p1_array_index_59081;
  reg [31:0] p1_array_index_59082;
  reg [31:0] p1_array_index_59084;
  reg [31:0] p1_array_index_59085;
  reg [31:0] p1_array_index_59089;
  reg [31:0] p1_array_index_59090;
  reg [31:0] p1_array_index_59092;
  reg [31:0] p1_array_index_59093;
  reg [31:0] p1_array_index_59097;
  reg [31:0] p1_array_index_59098;
  reg [31:0] p1_array_index_59100;
  reg [31:0] p1_array_index_59101;
  reg [31:0] p1_array_index_58978;
  reg [31:0] p1_array_index_58979;
  reg [31:0] p1_array_index_58984;
  reg [31:0] p1_array_index_58985;
  reg [31:0] p1_array_index_58992;
  reg [31:0] p1_array_index_58995;
  reg [31:0] p1_array_index_59000;
  reg [31:0] p1_array_index_59003;
  reg [31:0] p1_array_index_59008;
  reg [31:0] p1_array_index_59011;
  reg [31:0] p1_array_index_59016;
  reg [31:0] p1_array_index_59019;
  reg [31:0] p1_array_index_59024;
  reg [31:0] p1_array_index_59027;
  reg [31:0] p1_array_index_59032;
  reg [31:0] p1_array_index_59035;
  reg [31:0] p1_array_index_59040;
  reg [31:0] p1_array_index_59043;
  reg [31:0] p1_array_index_59048;
  reg [31:0] p1_array_index_59051;
  reg [31:0] p1_array_index_59056;
  reg [31:0] p1_array_index_59059;
  reg [31:0] p1_array_index_59064;
  reg [31:0] p1_array_index_59067;
  reg [31:0] p1_array_index_59072;
  reg [31:0] p1_array_index_59075;
  reg [31:0] p1_array_index_59080;
  reg [31:0] p1_array_index_59083;
  reg [31:0] p1_array_index_59088;
  reg [31:0] p1_array_index_59091;
  reg [31:0] p1_array_index_59096;
  reg [31:0] p1_array_index_59099;
  reg [31:0] p1_array_index_58976;
  reg [31:0] p1_array_index_58977;
  reg [31:0] p1_array_index_58991;
  reg [31:0] p1_array_index_58999;
  reg [31:0] p1_array_index_59007;
  reg [31:0] p1_array_index_59015;
  reg [31:0] p1_array_index_59023;
  reg [31:0] p1_array_index_59031;
  reg [31:0] p1_array_index_59039;
  reg [31:0] p1_array_index_59047;
  reg [31:0] p1_array_index_59055;
  reg [31:0] p1_array_index_59063;
  reg [31:0] p1_array_index_59071;
  reg [31:0] p1_array_index_59079;
  reg [31:0] p1_array_index_59087;
  reg [31:0] p1_array_index_59095;
  reg [31:0] p1_array_index_58974;
  reg [31:0] p1_array_index_58975;
  reg [31:0] p1_array_index_58990;
  reg [31:0] p1_array_index_58998;
  reg [31:0] p1_array_index_59006;
  reg [31:0] p1_array_index_59014;
  reg [31:0] p1_array_index_59022;
  reg [31:0] p1_array_index_59030;
  reg [31:0] p1_array_index_59038;
  reg [31:0] p1_array_index_59046;
  reg [31:0] p1_array_index_59054;
  reg [31:0] p1_array_index_59062;
  reg [31:0] p1_array_index_59070;
  reg [31:0] p1_array_index_59078;
  reg [31:0] p1_array_index_59086;
  reg [31:0] p1_array_index_59094;
  always_ff @ (posedge clk) begin
    p1_a <= p0_a;
    p1_b <= p0_b;
    p1_array_index_58980 <= p1_array_index_58980_comb;
    p1_array_index_58981 <= p1_array_index_58981_comb;
    p1_array_index_58982 <= p1_array_index_58982_comb;
    p1_array_index_58983 <= p1_array_index_58983_comb;
    p1_array_index_58986 <= p1_array_index_58986_comb;
    p1_array_index_58987 <= p1_array_index_58987_comb;
    p1_array_index_58988 <= p1_array_index_58988_comb;
    p1_array_index_58989 <= p1_array_index_58989_comb;
    p1_array_index_58993 <= p1_array_index_58993_comb;
    p1_array_index_58994 <= p1_array_index_58994_comb;
    p1_array_index_58996 <= p1_array_index_58996_comb;
    p1_array_index_58997 <= p1_array_index_58997_comb;
    p1_array_index_59001 <= p1_array_index_59001_comb;
    p1_array_index_59002 <= p1_array_index_59002_comb;
    p1_array_index_59004 <= p1_array_index_59004_comb;
    p1_array_index_59005 <= p1_array_index_59005_comb;
    p1_array_index_59009 <= p1_array_index_59009_comb;
    p1_array_index_59010 <= p1_array_index_59010_comb;
    p1_array_index_59012 <= p1_array_index_59012_comb;
    p1_array_index_59013 <= p1_array_index_59013_comb;
    p1_array_index_59017 <= p1_array_index_59017_comb;
    p1_array_index_59018 <= p1_array_index_59018_comb;
    p1_array_index_59020 <= p1_array_index_59020_comb;
    p1_array_index_59021 <= p1_array_index_59021_comb;
    p1_array_index_59025 <= p1_array_index_59025_comb;
    p1_array_index_59026 <= p1_array_index_59026_comb;
    p1_array_index_59028 <= p1_array_index_59028_comb;
    p1_array_index_59029 <= p1_array_index_59029_comb;
    p1_array_index_59033 <= p1_array_index_59033_comb;
    p1_array_index_59034 <= p1_array_index_59034_comb;
    p1_array_index_59036 <= p1_array_index_59036_comb;
    p1_array_index_59037 <= p1_array_index_59037_comb;
    p1_array_index_59041 <= p1_array_index_59041_comb;
    p1_array_index_59042 <= p1_array_index_59042_comb;
    p1_array_index_59044 <= p1_array_index_59044_comb;
    p1_array_index_59045 <= p1_array_index_59045_comb;
    p1_array_index_59049 <= p1_array_index_59049_comb;
    p1_array_index_59050 <= p1_array_index_59050_comb;
    p1_array_index_59052 <= p1_array_index_59052_comb;
    p1_array_index_59053 <= p1_array_index_59053_comb;
    p1_array_index_59057 <= p1_array_index_59057_comb;
    p1_array_index_59058 <= p1_array_index_59058_comb;
    p1_array_index_59060 <= p1_array_index_59060_comb;
    p1_array_index_59061 <= p1_array_index_59061_comb;
    p1_array_index_59065 <= p1_array_index_59065_comb;
    p1_array_index_59066 <= p1_array_index_59066_comb;
    p1_array_index_59068 <= p1_array_index_59068_comb;
    p1_array_index_59069 <= p1_array_index_59069_comb;
    p1_array_index_59073 <= p1_array_index_59073_comb;
    p1_array_index_59074 <= p1_array_index_59074_comb;
    p1_array_index_59076 <= p1_array_index_59076_comb;
    p1_array_index_59077 <= p1_array_index_59077_comb;
    p1_array_index_59081 <= p1_array_index_59081_comb;
    p1_array_index_59082 <= p1_array_index_59082_comb;
    p1_array_index_59084 <= p1_array_index_59084_comb;
    p1_array_index_59085 <= p1_array_index_59085_comb;
    p1_array_index_59089 <= p1_array_index_59089_comb;
    p1_array_index_59090 <= p1_array_index_59090_comb;
    p1_array_index_59092 <= p1_array_index_59092_comb;
    p1_array_index_59093 <= p1_array_index_59093_comb;
    p1_array_index_59097 <= p1_array_index_59097_comb;
    p1_array_index_59098 <= p1_array_index_59098_comb;
    p1_array_index_59100 <= p1_array_index_59100_comb;
    p1_array_index_59101 <= p1_array_index_59101_comb;
    p1_array_index_58978 <= p1_array_index_58978_comb;
    p1_array_index_58979 <= p1_array_index_58979_comb;
    p1_array_index_58984 <= p1_array_index_58984_comb;
    p1_array_index_58985 <= p1_array_index_58985_comb;
    p1_array_index_58992 <= p1_array_index_58992_comb;
    p1_array_index_58995 <= p1_array_index_58995_comb;
    p1_array_index_59000 <= p1_array_index_59000_comb;
    p1_array_index_59003 <= p1_array_index_59003_comb;
    p1_array_index_59008 <= p1_array_index_59008_comb;
    p1_array_index_59011 <= p1_array_index_59011_comb;
    p1_array_index_59016 <= p1_array_index_59016_comb;
    p1_array_index_59019 <= p1_array_index_59019_comb;
    p1_array_index_59024 <= p1_array_index_59024_comb;
    p1_array_index_59027 <= p1_array_index_59027_comb;
    p1_array_index_59032 <= p1_array_index_59032_comb;
    p1_array_index_59035 <= p1_array_index_59035_comb;
    p1_array_index_59040 <= p1_array_index_59040_comb;
    p1_array_index_59043 <= p1_array_index_59043_comb;
    p1_array_index_59048 <= p1_array_index_59048_comb;
    p1_array_index_59051 <= p1_array_index_59051_comb;
    p1_array_index_59056 <= p1_array_index_59056_comb;
    p1_array_index_59059 <= p1_array_index_59059_comb;
    p1_array_index_59064 <= p1_array_index_59064_comb;
    p1_array_index_59067 <= p1_array_index_59067_comb;
    p1_array_index_59072 <= p1_array_index_59072_comb;
    p1_array_index_59075 <= p1_array_index_59075_comb;
    p1_array_index_59080 <= p1_array_index_59080_comb;
    p1_array_index_59083 <= p1_array_index_59083_comb;
    p1_array_index_59088 <= p1_array_index_59088_comb;
    p1_array_index_59091 <= p1_array_index_59091_comb;
    p1_array_index_59096 <= p1_array_index_59096_comb;
    p1_array_index_59099 <= p1_array_index_59099_comb;
    p1_array_index_58976 <= p1_array_index_58976_comb;
    p1_array_index_58977 <= p1_array_index_58977_comb;
    p1_array_index_58991 <= p1_array_index_58991_comb;
    p1_array_index_58999 <= p1_array_index_58999_comb;
    p1_array_index_59007 <= p1_array_index_59007_comb;
    p1_array_index_59015 <= p1_array_index_59015_comb;
    p1_array_index_59023 <= p1_array_index_59023_comb;
    p1_array_index_59031 <= p1_array_index_59031_comb;
    p1_array_index_59039 <= p1_array_index_59039_comb;
    p1_array_index_59047 <= p1_array_index_59047_comb;
    p1_array_index_59055 <= p1_array_index_59055_comb;
    p1_array_index_59063 <= p1_array_index_59063_comb;
    p1_array_index_59071 <= p1_array_index_59071_comb;
    p1_array_index_59079 <= p1_array_index_59079_comb;
    p1_array_index_59087 <= p1_array_index_59087_comb;
    p1_array_index_59095 <= p1_array_index_59095_comb;
    p1_array_index_58974 <= p1_array_index_58974_comb;
    p1_array_index_58975 <= p1_array_index_58975_comb;
    p1_array_index_58990 <= p1_array_index_58990_comb;
    p1_array_index_58998 <= p1_array_index_58998_comb;
    p1_array_index_59006 <= p1_array_index_59006_comb;
    p1_array_index_59014 <= p1_array_index_59014_comb;
    p1_array_index_59022 <= p1_array_index_59022_comb;
    p1_array_index_59030 <= p1_array_index_59030_comb;
    p1_array_index_59038 <= p1_array_index_59038_comb;
    p1_array_index_59046 <= p1_array_index_59046_comb;
    p1_array_index_59054 <= p1_array_index_59054_comb;
    p1_array_index_59062 <= p1_array_index_59062_comb;
    p1_array_index_59070 <= p1_array_index_59070_comb;
    p1_array_index_59078 <= p1_array_index_59078_comb;
    p1_array_index_59086 <= p1_array_index_59086_comb;
    p1_array_index_59094 <= p1_array_index_59094_comb;
  end

  // ===== Pipe stage 2:
  wire [31:0] p2_smul_59866_comb;
  wire [31:0] p2_smul_59867_comb;
  wire [31:0] p2_smul_59868_comb;
  wire [31:0] p2_smul_59869_comb;
  wire [31:0] p2_smul_59870_comb;
  wire [31:0] p2_smul_59871_comb;
  wire [31:0] p2_smul_59872_comb;
  wire [31:0] p2_smul_59873_comb;
  wire [31:0] p2_smul_59858_comb;
  wire [31:0] p2_smul_59859_comb;
  wire [31:0] p2_smul_59860_comb;
  wire [31:0] p2_smul_59861_comb;
  wire [31:0] p2_smul_59862_comb;
  wire [31:0] p2_smul_59863_comb;
  wire [31:0] p2_smul_59864_comb;
  wire [31:0] p2_smul_59865_comb;
  wire [31:0] p2_smul_59850_comb;
  wire [31:0] p2_smul_59851_comb;
  wire [31:0] p2_smul_59852_comb;
  wire [31:0] p2_smul_59853_comb;
  wire [31:0] p2_smul_59854_comb;
  wire [31:0] p2_smul_59855_comb;
  wire [31:0] p2_smul_59856_comb;
  wire [31:0] p2_smul_59857_comb;
  wire [31:0] p2_smul_59842_comb;
  wire [31:0] p2_smul_59843_comb;
  wire [31:0] p2_smul_59844_comb;
  wire [31:0] p2_smul_59845_comb;
  wire [31:0] p2_smul_59846_comb;
  wire [31:0] p2_smul_59847_comb;
  wire [31:0] p2_smul_59848_comb;
  wire [31:0] p2_smul_59849_comb;
  wire [31:0] p2_smul_59834_comb;
  wire [31:0] p2_smul_59835_comb;
  wire [31:0] p2_smul_59836_comb;
  wire [31:0] p2_smul_59837_comb;
  wire [31:0] p2_smul_59838_comb;
  wire [31:0] p2_smul_59839_comb;
  wire [31:0] p2_smul_59840_comb;
  wire [31:0] p2_smul_59841_comb;
  wire [31:0] p2_smul_59826_comb;
  wire [31:0] p2_smul_59827_comb;
  wire [31:0] p2_smul_59828_comb;
  wire [31:0] p2_smul_59829_comb;
  wire [31:0] p2_smul_59830_comb;
  wire [31:0] p2_smul_59831_comb;
  wire [31:0] p2_smul_59832_comb;
  wire [31:0] p2_smul_59833_comb;
  wire [31:0] p2_smul_59818_comb;
  wire [31:0] p2_smul_59819_comb;
  wire [31:0] p2_smul_59820_comb;
  wire [31:0] p2_smul_59821_comb;
  wire [31:0] p2_smul_59822_comb;
  wire [31:0] p2_smul_59823_comb;
  wire [31:0] p2_smul_59824_comb;
  wire [31:0] p2_smul_59825_comb;
  wire [31:0] p2_smul_59810_comb;
  wire [31:0] p2_smul_59811_comb;
  wire [31:0] p2_smul_59812_comb;
  wire [31:0] p2_smul_59813_comb;
  wire [31:0] p2_smul_59814_comb;
  wire [31:0] p2_smul_59815_comb;
  wire [31:0] p2_smul_59816_comb;
  wire [31:0] p2_smul_59817_comb;
  wire [31:0] p2_smul_59802_comb;
  wire [31:0] p2_smul_59803_comb;
  wire [31:0] p2_smul_59804_comb;
  wire [31:0] p2_smul_59805_comb;
  wire [31:0] p2_smul_59806_comb;
  wire [31:0] p2_smul_59807_comb;
  wire [31:0] p2_smul_59808_comb;
  wire [31:0] p2_smul_59809_comb;
  wire [31:0] p2_smul_59794_comb;
  wire [31:0] p2_smul_59795_comb;
  wire [31:0] p2_smul_59796_comb;
  wire [31:0] p2_smul_59797_comb;
  wire [31:0] p2_smul_59798_comb;
  wire [31:0] p2_smul_59799_comb;
  wire [31:0] p2_smul_59800_comb;
  wire [31:0] p2_smul_59801_comb;
  wire [31:0] p2_smul_59786_comb;
  wire [31:0] p2_smul_59787_comb;
  wire [31:0] p2_smul_59788_comb;
  wire [31:0] p2_smul_59789_comb;
  wire [31:0] p2_smul_59790_comb;
  wire [31:0] p2_smul_59791_comb;
  wire [31:0] p2_smul_59792_comb;
  wire [31:0] p2_smul_59793_comb;
  wire [31:0] p2_smul_59778_comb;
  wire [31:0] p2_smul_59779_comb;
  wire [31:0] p2_smul_59780_comb;
  wire [31:0] p2_smul_59781_comb;
  wire [31:0] p2_smul_59782_comb;
  wire [31:0] p2_smul_59783_comb;
  wire [31:0] p2_smul_59784_comb;
  wire [31:0] p2_smul_59785_comb;
  wire [31:0] p2_smul_59770_comb;
  wire [31:0] p2_smul_59771_comb;
  wire [31:0] p2_smul_59772_comb;
  wire [31:0] p2_smul_59773_comb;
  wire [31:0] p2_smul_59774_comb;
  wire [31:0] p2_smul_59775_comb;
  wire [31:0] p2_smul_59776_comb;
  wire [31:0] p2_smul_59777_comb;
  wire [31:0] p2_smul_59762_comb;
  wire [31:0] p2_smul_59763_comb;
  wire [31:0] p2_smul_59764_comb;
  wire [31:0] p2_smul_59765_comb;
  wire [31:0] p2_smul_59766_comb;
  wire [31:0] p2_smul_59767_comb;
  wire [31:0] p2_smul_59768_comb;
  wire [31:0] p2_smul_59769_comb;
  wire [31:0] p2_smul_59754_comb;
  wire [31:0] p2_smul_59755_comb;
  wire [31:0] p2_smul_59756_comb;
  wire [31:0] p2_smul_59757_comb;
  wire [31:0] p2_smul_59758_comb;
  wire [31:0] p2_smul_59759_comb;
  wire [31:0] p2_smul_59760_comb;
  wire [31:0] p2_smul_59761_comb;
  wire [31:0] p2_smul_59746_comb;
  wire [31:0] p2_smul_59747_comb;
  wire [31:0] p2_smul_59748_comb;
  wire [31:0] p2_smul_59749_comb;
  wire [31:0] p2_smul_59750_comb;
  wire [31:0] p2_smul_59751_comb;
  wire [31:0] p2_smul_59752_comb;
  wire [31:0] p2_smul_59753_comb;
  wire [31:0] p2_smul_59738_comb;
  wire [31:0] p2_smul_59739_comb;
  wire [31:0] p2_smul_59740_comb;
  wire [31:0] p2_smul_59741_comb;
  wire [31:0] p2_smul_59742_comb;
  wire [31:0] p2_smul_59743_comb;
  wire [31:0] p2_smul_59744_comb;
  wire [31:0] p2_smul_59745_comb;
  wire [31:0] p2_smul_59730_comb;
  wire [31:0] p2_smul_59731_comb;
  wire [31:0] p2_smul_59732_comb;
  wire [31:0] p2_smul_59733_comb;
  wire [31:0] p2_smul_59734_comb;
  wire [31:0] p2_smul_59735_comb;
  wire [31:0] p2_smul_59736_comb;
  wire [31:0] p2_smul_59737_comb;
  wire [31:0] p2_smul_59722_comb;
  wire [31:0] p2_smul_59723_comb;
  wire [31:0] p2_smul_59724_comb;
  wire [31:0] p2_smul_59725_comb;
  wire [31:0] p2_smul_59726_comb;
  wire [31:0] p2_smul_59727_comb;
  wire [31:0] p2_smul_59728_comb;
  wire [31:0] p2_smul_59729_comb;
  wire [31:0] p2_smul_59714_comb;
  wire [31:0] p2_smul_59715_comb;
  wire [31:0] p2_smul_59716_comb;
  wire [31:0] p2_smul_59717_comb;
  wire [31:0] p2_smul_59718_comb;
  wire [31:0] p2_smul_59719_comb;
  wire [31:0] p2_smul_59720_comb;
  wire [31:0] p2_smul_59721_comb;
  wire [31:0] p2_smul_59706_comb;
  wire [31:0] p2_smul_59707_comb;
  wire [31:0] p2_smul_59708_comb;
  wire [31:0] p2_smul_59709_comb;
  wire [31:0] p2_smul_59710_comb;
  wire [31:0] p2_smul_59711_comb;
  wire [31:0] p2_smul_59712_comb;
  wire [31:0] p2_smul_59713_comb;
  wire [31:0] p2_smul_59698_comb;
  wire [31:0] p2_smul_59699_comb;
  wire [31:0] p2_smul_59700_comb;
  wire [31:0] p2_smul_59701_comb;
  wire [31:0] p2_smul_59702_comb;
  wire [31:0] p2_smul_59703_comb;
  wire [31:0] p2_smul_59704_comb;
  wire [31:0] p2_smul_59705_comb;
  wire [31:0] p2_smul_59690_comb;
  wire [31:0] p2_smul_59691_comb;
  wire [31:0] p2_smul_59692_comb;
  wire [31:0] p2_smul_59693_comb;
  wire [31:0] p2_smul_59694_comb;
  wire [31:0] p2_smul_59695_comb;
  wire [31:0] p2_smul_59696_comb;
  wire [31:0] p2_smul_59697_comb;
  wire [31:0] p2_smul_59682_comb;
  wire [31:0] p2_smul_59683_comb;
  wire [31:0] p2_smul_59684_comb;
  wire [31:0] p2_smul_59685_comb;
  wire [31:0] p2_smul_59686_comb;
  wire [31:0] p2_smul_59687_comb;
  wire [31:0] p2_smul_59688_comb;
  wire [31:0] p2_smul_59689_comb;
  wire [31:0] p2_smul_59674_comb;
  wire [31:0] p2_smul_59675_comb;
  wire [31:0] p2_smul_59676_comb;
  wire [31:0] p2_smul_59677_comb;
  wire [31:0] p2_smul_59678_comb;
  wire [31:0] p2_smul_59679_comb;
  wire [31:0] p2_smul_59680_comb;
  wire [31:0] p2_smul_59681_comb;
  wire [31:0] p2_smul_59666_comb;
  wire [31:0] p2_smul_59667_comb;
  wire [31:0] p2_smul_59668_comb;
  wire [31:0] p2_smul_59669_comb;
  wire [31:0] p2_smul_59670_comb;
  wire [31:0] p2_smul_59671_comb;
  wire [31:0] p2_smul_59672_comb;
  wire [31:0] p2_smul_59673_comb;
  wire [31:0] p2_smul_59658_comb;
  wire [31:0] p2_smul_59659_comb;
  wire [31:0] p2_smul_59660_comb;
  wire [31:0] p2_smul_59661_comb;
  wire [31:0] p2_smul_59662_comb;
  wire [31:0] p2_smul_59663_comb;
  wire [31:0] p2_smul_59664_comb;
  wire [31:0] p2_smul_59665_comb;
  wire [31:0] p2_smul_59650_comb;
  wire [31:0] p2_smul_59651_comb;
  wire [31:0] p2_smul_59652_comb;
  wire [31:0] p2_smul_59653_comb;
  wire [31:0] p2_smul_59654_comb;
  wire [31:0] p2_smul_59655_comb;
  wire [31:0] p2_smul_59656_comb;
  wire [31:0] p2_smul_59657_comb;
  wire [31:0] p2_smul_59642_comb;
  wire [31:0] p2_smul_59643_comb;
  wire [31:0] p2_smul_59644_comb;
  wire [31:0] p2_smul_59645_comb;
  wire [31:0] p2_smul_59646_comb;
  wire [31:0] p2_smul_59647_comb;
  wire [31:0] p2_smul_59648_comb;
  wire [31:0] p2_smul_59649_comb;
  wire [31:0] p2_smul_59634_comb;
  wire [31:0] p2_smul_59635_comb;
  wire [31:0] p2_smul_59636_comb;
  wire [31:0] p2_smul_59637_comb;
  wire [31:0] p2_smul_59638_comb;
  wire [31:0] p2_smul_59639_comb;
  wire [31:0] p2_smul_59640_comb;
  wire [31:0] p2_smul_59641_comb;
  wire [31:0] p2_smul_59626_comb;
  wire [31:0] p2_smul_59627_comb;
  wire [31:0] p2_smul_59628_comb;
  wire [31:0] p2_smul_59629_comb;
  wire [31:0] p2_smul_59630_comb;
  wire [31:0] p2_smul_59631_comb;
  wire [31:0] p2_smul_59632_comb;
  wire [31:0] p2_smul_59633_comb;
  wire [31:0] p2_smul_59618_comb;
  wire [31:0] p2_smul_59619_comb;
  wire [31:0] p2_smul_59620_comb;
  wire [31:0] p2_smul_59621_comb;
  wire [31:0] p2_smul_59622_comb;
  wire [31:0] p2_smul_59623_comb;
  wire [31:0] p2_smul_59624_comb;
  wire [31:0] p2_smul_59625_comb;
  wire [31:0] p2_smul_59610_comb;
  wire [31:0] p2_smul_59611_comb;
  wire [31:0] p2_smul_59612_comb;
  wire [31:0] p2_smul_59613_comb;
  wire [31:0] p2_smul_59614_comb;
  wire [31:0] p2_smul_59615_comb;
  wire [31:0] p2_smul_59616_comb;
  wire [31:0] p2_smul_59617_comb;
  wire [31:0] p2_smul_59602_comb;
  wire [31:0] p2_smul_59603_comb;
  wire [31:0] p2_smul_59604_comb;
  wire [31:0] p2_smul_59605_comb;
  wire [31:0] p2_smul_59606_comb;
  wire [31:0] p2_smul_59607_comb;
  wire [31:0] p2_smul_59608_comb;
  wire [31:0] p2_smul_59609_comb;
  wire [31:0] p2_smul_59594_comb;
  wire [31:0] p2_smul_59595_comb;
  wire [31:0] p2_smul_59596_comb;
  wire [31:0] p2_smul_59597_comb;
  wire [31:0] p2_smul_59598_comb;
  wire [31:0] p2_smul_59599_comb;
  wire [31:0] p2_smul_59600_comb;
  wire [31:0] p2_smul_59601_comb;
  wire [31:0] p2_smul_59586_comb;
  wire [31:0] p2_smul_59587_comb;
  wire [31:0] p2_smul_59588_comb;
  wire [31:0] p2_smul_59589_comb;
  wire [31:0] p2_smul_59590_comb;
  wire [31:0] p2_smul_59591_comb;
  wire [31:0] p2_smul_59592_comb;
  wire [31:0] p2_smul_59593_comb;
  wire [31:0] p2_smul_59578_comb;
  wire [31:0] p2_smul_59579_comb;
  wire [31:0] p2_smul_59580_comb;
  wire [31:0] p2_smul_59581_comb;
  wire [31:0] p2_smul_59582_comb;
  wire [31:0] p2_smul_59583_comb;
  wire [31:0] p2_smul_59584_comb;
  wire [31:0] p2_smul_59585_comb;
  wire [31:0] p2_smul_59570_comb;
  wire [31:0] p2_smul_59571_comb;
  wire [31:0] p2_smul_59572_comb;
  wire [31:0] p2_smul_59573_comb;
  wire [31:0] p2_smul_59574_comb;
  wire [31:0] p2_smul_59575_comb;
  wire [31:0] p2_smul_59576_comb;
  wire [31:0] p2_smul_59577_comb;
  wire [31:0] p2_smul_59562_comb;
  wire [31:0] p2_smul_59563_comb;
  wire [31:0] p2_smul_59564_comb;
  wire [31:0] p2_smul_59565_comb;
  wire [31:0] p2_smul_59566_comb;
  wire [31:0] p2_smul_59567_comb;
  wire [31:0] p2_smul_59568_comb;
  wire [31:0] p2_smul_59569_comb;
  wire [31:0] p2_smul_59554_comb;
  wire [31:0] p2_smul_59555_comb;
  wire [31:0] p2_smul_59556_comb;
  wire [31:0] p2_smul_59557_comb;
  wire [31:0] p2_smul_59558_comb;
  wire [31:0] p2_smul_59559_comb;
  wire [31:0] p2_smul_59560_comb;
  wire [31:0] p2_smul_59561_comb;
  wire [31:0] p2_smul_59546_comb;
  wire [31:0] p2_smul_59547_comb;
  wire [31:0] p2_smul_59548_comb;
  wire [31:0] p2_smul_59549_comb;
  wire [31:0] p2_smul_59550_comb;
  wire [31:0] p2_smul_59551_comb;
  wire [31:0] p2_smul_59552_comb;
  wire [31:0] p2_smul_59553_comb;
  wire [31:0] p2_smul_59538_comb;
  wire [31:0] p2_smul_59539_comb;
  wire [31:0] p2_smul_59540_comb;
  wire [31:0] p2_smul_59541_comb;
  wire [31:0] p2_smul_59542_comb;
  wire [31:0] p2_smul_59543_comb;
  wire [31:0] p2_smul_59544_comb;
  wire [31:0] p2_smul_59545_comb;
  wire [31:0] p2_smul_59530_comb;
  wire [31:0] p2_smul_59531_comb;
  wire [31:0] p2_smul_59532_comb;
  wire [31:0] p2_smul_59533_comb;
  wire [31:0] p2_smul_59534_comb;
  wire [31:0] p2_smul_59535_comb;
  wire [31:0] p2_smul_59536_comb;
  wire [31:0] p2_smul_59537_comb;
  wire [31:0] p2_smul_59522_comb;
  wire [31:0] p2_smul_59523_comb;
  wire [31:0] p2_smul_59524_comb;
  wire [31:0] p2_smul_59525_comb;
  wire [31:0] p2_smul_59526_comb;
  wire [31:0] p2_smul_59527_comb;
  wire [31:0] p2_smul_59528_comb;
  wire [31:0] p2_smul_59529_comb;
  wire [31:0] p2_smul_59514_comb;
  wire [31:0] p2_smul_59515_comb;
  wire [31:0] p2_smul_59516_comb;
  wire [31:0] p2_smul_59517_comb;
  wire [31:0] p2_smul_59518_comb;
  wire [31:0] p2_smul_59519_comb;
  wire [31:0] p2_smul_59520_comb;
  wire [31:0] p2_smul_59521_comb;
  wire [31:0] p2_smul_59506_comb;
  wire [31:0] p2_smul_59507_comb;
  wire [31:0] p2_smul_59508_comb;
  wire [31:0] p2_smul_59509_comb;
  wire [31:0] p2_smul_59510_comb;
  wire [31:0] p2_smul_59511_comb;
  wire [31:0] p2_smul_59512_comb;
  wire [31:0] p2_smul_59513_comb;
  wire [31:0] p2_smul_59498_comb;
  wire [31:0] p2_smul_59499_comb;
  wire [31:0] p2_smul_59500_comb;
  wire [31:0] p2_smul_59501_comb;
  wire [31:0] p2_smul_59502_comb;
  wire [31:0] p2_smul_59503_comb;
  wire [31:0] p2_smul_59504_comb;
  wire [31:0] p2_smul_59505_comb;
  wire [31:0] p2_smul_59490_comb;
  wire [31:0] p2_smul_59491_comb;
  wire [31:0] p2_smul_59492_comb;
  wire [31:0] p2_smul_59493_comb;
  wire [31:0] p2_smul_59494_comb;
  wire [31:0] p2_smul_59495_comb;
  wire [31:0] p2_smul_59496_comb;
  wire [31:0] p2_smul_59497_comb;
  wire [31:0] p2_smul_59482_comb;
  wire [31:0] p2_smul_59483_comb;
  wire [31:0] p2_smul_59484_comb;
  wire [31:0] p2_smul_59485_comb;
  wire [31:0] p2_smul_59486_comb;
  wire [31:0] p2_smul_59487_comb;
  wire [31:0] p2_smul_59488_comb;
  wire [31:0] p2_smul_59489_comb;
  wire [31:0] p2_smul_59474_comb;
  wire [31:0] p2_smul_59475_comb;
  wire [31:0] p2_smul_59476_comb;
  wire [31:0] p2_smul_59477_comb;
  wire [31:0] p2_smul_59478_comb;
  wire [31:0] p2_smul_59479_comb;
  wire [31:0] p2_smul_59480_comb;
  wire [31:0] p2_smul_59481_comb;
  wire [31:0] p2_smul_59466_comb;
  wire [31:0] p2_smul_59467_comb;
  wire [31:0] p2_smul_59468_comb;
  wire [31:0] p2_smul_59469_comb;
  wire [31:0] p2_smul_59470_comb;
  wire [31:0] p2_smul_59471_comb;
  wire [31:0] p2_smul_59472_comb;
  wire [31:0] p2_smul_59473_comb;
  wire [31:0] p2_smul_59458_comb;
  wire [31:0] p2_smul_59459_comb;
  wire [31:0] p2_smul_59460_comb;
  wire [31:0] p2_smul_59461_comb;
  wire [31:0] p2_smul_59462_comb;
  wire [31:0] p2_smul_59463_comb;
  wire [31:0] p2_smul_59464_comb;
  wire [31:0] p2_smul_59465_comb;
  wire [31:0] p2_smul_59450_comb;
  wire [31:0] p2_smul_59451_comb;
  wire [31:0] p2_smul_59452_comb;
  wire [31:0] p2_smul_59453_comb;
  wire [31:0] p2_smul_59454_comb;
  wire [31:0] p2_smul_59455_comb;
  wire [31:0] p2_smul_59456_comb;
  wire [31:0] p2_smul_59457_comb;
  wire [31:0] p2_smul_59442_comb;
  wire [31:0] p2_smul_59443_comb;
  wire [31:0] p2_smul_59444_comb;
  wire [31:0] p2_smul_59445_comb;
  wire [31:0] p2_smul_59446_comb;
  wire [31:0] p2_smul_59447_comb;
  wire [31:0] p2_smul_59448_comb;
  wire [31:0] p2_smul_59449_comb;
  wire [31:0] p2_smul_59434_comb;
  wire [31:0] p2_smul_59435_comb;
  wire [31:0] p2_smul_59436_comb;
  wire [31:0] p2_smul_59437_comb;
  wire [31:0] p2_smul_59438_comb;
  wire [31:0] p2_smul_59439_comb;
  wire [31:0] p2_smul_59440_comb;
  wire [31:0] p2_smul_59441_comb;
  wire [31:0] p2_smul_59426_comb;
  wire [31:0] p2_smul_59427_comb;
  wire [31:0] p2_smul_59428_comb;
  wire [31:0] p2_smul_59429_comb;
  wire [31:0] p2_smul_59430_comb;
  wire [31:0] p2_smul_59431_comb;
  wire [31:0] p2_smul_59432_comb;
  wire [31:0] p2_smul_59433_comb;
  wire [31:0] p2_smul_59418_comb;
  wire [31:0] p2_smul_59419_comb;
  wire [31:0] p2_smul_59420_comb;
  wire [31:0] p2_smul_59421_comb;
  wire [31:0] p2_smul_59422_comb;
  wire [31:0] p2_smul_59423_comb;
  wire [31:0] p2_smul_59424_comb;
  wire [31:0] p2_smul_59425_comb;
  wire [31:0] p2_smul_59410_comb;
  wire [31:0] p2_smul_59411_comb;
  wire [31:0] p2_smul_59412_comb;
  wire [31:0] p2_smul_59413_comb;
  wire [31:0] p2_smul_59414_comb;
  wire [31:0] p2_smul_59415_comb;
  wire [31:0] p2_smul_59416_comb;
  wire [31:0] p2_smul_59417_comb;
  wire [31:0] p2_smul_59402_comb;
  wire [31:0] p2_smul_59403_comb;
  wire [31:0] p2_smul_59404_comb;
  wire [31:0] p2_smul_59405_comb;
  wire [31:0] p2_smul_59406_comb;
  wire [31:0] p2_smul_59407_comb;
  wire [31:0] p2_smul_59408_comb;
  wire [31:0] p2_smul_59409_comb;
  wire [31:0] p2_smul_59394_comb;
  wire [31:0] p2_smul_59395_comb;
  wire [31:0] p2_smul_59396_comb;
  wire [31:0] p2_smul_59397_comb;
  wire [31:0] p2_smul_59398_comb;
  wire [31:0] p2_smul_59399_comb;
  wire [31:0] p2_smul_59400_comb;
  wire [31:0] p2_smul_59401_comb;
  wire [31:0] p2_smul_59386_comb;
  wire [31:0] p2_smul_59387_comb;
  wire [31:0] p2_smul_59388_comb;
  wire [31:0] p2_smul_59389_comb;
  wire [31:0] p2_smul_59390_comb;
  wire [31:0] p2_smul_59391_comb;
  wire [31:0] p2_smul_59392_comb;
  wire [31:0] p2_smul_59393_comb;
  wire [31:0] p2_smul_59378_comb;
  wire [31:0] p2_smul_59379_comb;
  wire [31:0] p2_smul_59380_comb;
  wire [31:0] p2_smul_59381_comb;
  wire [31:0] p2_smul_59382_comb;
  wire [31:0] p2_smul_59383_comb;
  wire [31:0] p2_smul_59384_comb;
  wire [31:0] p2_smul_59385_comb;
  wire [31:0] p2_smul_59370_comb;
  wire [31:0] p2_smul_59371_comb;
  wire [31:0] p2_smul_59372_comb;
  wire [31:0] p2_smul_59373_comb;
  wire [31:0] p2_smul_59374_comb;
  wire [31:0] p2_smul_59375_comb;
  wire [31:0] p2_smul_59376_comb;
  wire [31:0] p2_smul_59377_comb;
  wire [31:0] p2_smul_59362_comb;
  wire [31:0] p2_smul_59363_comb;
  wire [31:0] p2_smul_59364_comb;
  wire [31:0] p2_smul_59365_comb;
  wire [31:0] p2_smul_59366_comb;
  wire [31:0] p2_smul_59367_comb;
  wire [31:0] p2_smul_59368_comb;
  wire [31:0] p2_smul_59369_comb;
  wire [31:0] p2_add_60126_comb;
  wire [31:0] p2_add_60127_comb;
  wire [31:0] p2_add_60128_comb;
  wire [31:0] p2_add_60129_comb;
  wire [31:0] p2_add_60122_comb;
  wire [31:0] p2_add_60123_comb;
  wire [31:0] p2_add_60124_comb;
  wire [31:0] p2_add_60125_comb;
  wire [31:0] p2_add_60118_comb;
  wire [31:0] p2_add_60119_comb;
  wire [31:0] p2_add_60120_comb;
  wire [31:0] p2_add_60121_comb;
  wire [31:0] p2_add_60114_comb;
  wire [31:0] p2_add_60115_comb;
  wire [31:0] p2_add_60116_comb;
  wire [31:0] p2_add_60117_comb;
  wire [31:0] p2_add_60110_comb;
  wire [31:0] p2_add_60111_comb;
  wire [31:0] p2_add_60112_comb;
  wire [31:0] p2_add_60113_comb;
  wire [31:0] p2_add_60106_comb;
  wire [31:0] p2_add_60107_comb;
  wire [31:0] p2_add_60108_comb;
  wire [31:0] p2_add_60109_comb;
  wire [31:0] p2_add_60102_comb;
  wire [31:0] p2_add_60103_comb;
  wire [31:0] p2_add_60104_comb;
  wire [31:0] p2_add_60105_comb;
  wire [31:0] p2_add_60098_comb;
  wire [31:0] p2_add_60099_comb;
  wire [31:0] p2_add_60100_comb;
  wire [31:0] p2_add_60101_comb;
  wire [31:0] p2_add_60094_comb;
  wire [31:0] p2_add_60095_comb;
  wire [31:0] p2_add_60096_comb;
  wire [31:0] p2_add_60097_comb;
  wire [31:0] p2_add_60090_comb;
  wire [31:0] p2_add_60091_comb;
  wire [31:0] p2_add_60092_comb;
  wire [31:0] p2_add_60093_comb;
  wire [31:0] p2_add_60086_comb;
  wire [31:0] p2_add_60087_comb;
  wire [31:0] p2_add_60088_comb;
  wire [31:0] p2_add_60089_comb;
  wire [31:0] p2_add_60082_comb;
  wire [31:0] p2_add_60083_comb;
  wire [31:0] p2_add_60084_comb;
  wire [31:0] p2_add_60085_comb;
  wire [31:0] p2_add_60078_comb;
  wire [31:0] p2_add_60079_comb;
  wire [31:0] p2_add_60080_comb;
  wire [31:0] p2_add_60081_comb;
  wire [31:0] p2_add_60074_comb;
  wire [31:0] p2_add_60075_comb;
  wire [31:0] p2_add_60076_comb;
  wire [31:0] p2_add_60077_comb;
  wire [31:0] p2_add_60070_comb;
  wire [31:0] p2_add_60071_comb;
  wire [31:0] p2_add_60072_comb;
  wire [31:0] p2_add_60073_comb;
  wire [31:0] p2_add_60066_comb;
  wire [31:0] p2_add_60067_comb;
  wire [31:0] p2_add_60068_comb;
  wire [31:0] p2_add_60069_comb;
  wire [31:0] p2_add_60062_comb;
  wire [31:0] p2_add_60063_comb;
  wire [31:0] p2_add_60064_comb;
  wire [31:0] p2_add_60065_comb;
  wire [31:0] p2_add_60058_comb;
  wire [31:0] p2_add_60059_comb;
  wire [31:0] p2_add_60060_comb;
  wire [31:0] p2_add_60061_comb;
  wire [31:0] p2_add_60054_comb;
  wire [31:0] p2_add_60055_comb;
  wire [31:0] p2_add_60056_comb;
  wire [31:0] p2_add_60057_comb;
  wire [31:0] p2_add_60050_comb;
  wire [31:0] p2_add_60051_comb;
  wire [31:0] p2_add_60052_comb;
  wire [31:0] p2_add_60053_comb;
  wire [31:0] p2_add_60046_comb;
  wire [31:0] p2_add_60047_comb;
  wire [31:0] p2_add_60048_comb;
  wire [31:0] p2_add_60049_comb;
  wire [31:0] p2_add_60042_comb;
  wire [31:0] p2_add_60043_comb;
  wire [31:0] p2_add_60044_comb;
  wire [31:0] p2_add_60045_comb;
  wire [31:0] p2_add_60038_comb;
  wire [31:0] p2_add_60039_comb;
  wire [31:0] p2_add_60040_comb;
  wire [31:0] p2_add_60041_comb;
  wire [31:0] p2_add_60034_comb;
  wire [31:0] p2_add_60035_comb;
  wire [31:0] p2_add_60036_comb;
  wire [31:0] p2_add_60037_comb;
  wire [31:0] p2_add_60030_comb;
  wire [31:0] p2_add_60031_comb;
  wire [31:0] p2_add_60032_comb;
  wire [31:0] p2_add_60033_comb;
  wire [31:0] p2_add_60026_comb;
  wire [31:0] p2_add_60027_comb;
  wire [31:0] p2_add_60028_comb;
  wire [31:0] p2_add_60029_comb;
  wire [31:0] p2_add_60022_comb;
  wire [31:0] p2_add_60023_comb;
  wire [31:0] p2_add_60024_comb;
  wire [31:0] p2_add_60025_comb;
  wire [31:0] p2_add_60018_comb;
  wire [31:0] p2_add_60019_comb;
  wire [31:0] p2_add_60020_comb;
  wire [31:0] p2_add_60021_comb;
  wire [31:0] p2_add_60014_comb;
  wire [31:0] p2_add_60015_comb;
  wire [31:0] p2_add_60016_comb;
  wire [31:0] p2_add_60017_comb;
  wire [31:0] p2_add_60010_comb;
  wire [31:0] p2_add_60011_comb;
  wire [31:0] p2_add_60012_comb;
  wire [31:0] p2_add_60013_comb;
  wire [31:0] p2_add_60006_comb;
  wire [31:0] p2_add_60007_comb;
  wire [31:0] p2_add_60008_comb;
  wire [31:0] p2_add_60009_comb;
  wire [31:0] p2_add_60002_comb;
  wire [31:0] p2_add_60003_comb;
  wire [31:0] p2_add_60004_comb;
  wire [31:0] p2_add_60005_comb;
  wire [31:0] p2_add_59998_comb;
  wire [31:0] p2_add_59999_comb;
  wire [31:0] p2_add_60000_comb;
  wire [31:0] p2_add_60001_comb;
  wire [31:0] p2_add_59994_comb;
  wire [31:0] p2_add_59995_comb;
  wire [31:0] p2_add_59996_comb;
  wire [31:0] p2_add_59997_comb;
  wire [31:0] p2_add_59990_comb;
  wire [31:0] p2_add_59991_comb;
  wire [31:0] p2_add_59992_comb;
  wire [31:0] p2_add_59993_comb;
  wire [31:0] p2_add_59986_comb;
  wire [31:0] p2_add_59987_comb;
  wire [31:0] p2_add_59988_comb;
  wire [31:0] p2_add_59989_comb;
  wire [31:0] p2_add_59982_comb;
  wire [31:0] p2_add_59983_comb;
  wire [31:0] p2_add_59984_comb;
  wire [31:0] p2_add_59985_comb;
  wire [31:0] p2_add_59978_comb;
  wire [31:0] p2_add_59979_comb;
  wire [31:0] p2_add_59980_comb;
  wire [31:0] p2_add_59981_comb;
  wire [31:0] p2_add_59974_comb;
  wire [31:0] p2_add_59975_comb;
  wire [31:0] p2_add_59976_comb;
  wire [31:0] p2_add_59977_comb;
  wire [31:0] p2_add_59970_comb;
  wire [31:0] p2_add_59971_comb;
  wire [31:0] p2_add_59972_comb;
  wire [31:0] p2_add_59973_comb;
  wire [31:0] p2_add_59966_comb;
  wire [31:0] p2_add_59967_comb;
  wire [31:0] p2_add_59968_comb;
  wire [31:0] p2_add_59969_comb;
  wire [31:0] p2_add_59962_comb;
  wire [31:0] p2_add_59963_comb;
  wire [31:0] p2_add_59964_comb;
  wire [31:0] p2_add_59965_comb;
  wire [31:0] p2_add_59958_comb;
  wire [31:0] p2_add_59959_comb;
  wire [31:0] p2_add_59960_comb;
  wire [31:0] p2_add_59961_comb;
  wire [31:0] p2_add_59954_comb;
  wire [31:0] p2_add_59955_comb;
  wire [31:0] p2_add_59956_comb;
  wire [31:0] p2_add_59957_comb;
  wire [31:0] p2_add_59950_comb;
  wire [31:0] p2_add_59951_comb;
  wire [31:0] p2_add_59952_comb;
  wire [31:0] p2_add_59953_comb;
  wire [31:0] p2_add_59946_comb;
  wire [31:0] p2_add_59947_comb;
  wire [31:0] p2_add_59948_comb;
  wire [31:0] p2_add_59949_comb;
  wire [31:0] p2_add_59942_comb;
  wire [31:0] p2_add_59943_comb;
  wire [31:0] p2_add_59944_comb;
  wire [31:0] p2_add_59945_comb;
  wire [31:0] p2_add_59938_comb;
  wire [31:0] p2_add_59939_comb;
  wire [31:0] p2_add_59940_comb;
  wire [31:0] p2_add_59941_comb;
  wire [31:0] p2_add_59934_comb;
  wire [31:0] p2_add_59935_comb;
  wire [31:0] p2_add_59936_comb;
  wire [31:0] p2_add_59937_comb;
  wire [31:0] p2_add_59930_comb;
  wire [31:0] p2_add_59931_comb;
  wire [31:0] p2_add_59932_comb;
  wire [31:0] p2_add_59933_comb;
  wire [31:0] p2_add_59926_comb;
  wire [31:0] p2_add_59927_comb;
  wire [31:0] p2_add_59928_comb;
  wire [31:0] p2_add_59929_comb;
  wire [31:0] p2_add_59922_comb;
  wire [31:0] p2_add_59923_comb;
  wire [31:0] p2_add_59924_comb;
  wire [31:0] p2_add_59925_comb;
  wire [31:0] p2_add_59918_comb;
  wire [31:0] p2_add_59919_comb;
  wire [31:0] p2_add_59920_comb;
  wire [31:0] p2_add_59921_comb;
  wire [31:0] p2_add_59914_comb;
  wire [31:0] p2_add_59915_comb;
  wire [31:0] p2_add_59916_comb;
  wire [31:0] p2_add_59917_comb;
  wire [31:0] p2_add_59910_comb;
  wire [31:0] p2_add_59911_comb;
  wire [31:0] p2_add_59912_comb;
  wire [31:0] p2_add_59913_comb;
  wire [31:0] p2_add_59906_comb;
  wire [31:0] p2_add_59907_comb;
  wire [31:0] p2_add_59908_comb;
  wire [31:0] p2_add_59909_comb;
  wire [31:0] p2_add_59902_comb;
  wire [31:0] p2_add_59903_comb;
  wire [31:0] p2_add_59904_comb;
  wire [31:0] p2_add_59905_comb;
  wire [31:0] p2_add_59898_comb;
  wire [31:0] p2_add_59899_comb;
  wire [31:0] p2_add_59900_comb;
  wire [31:0] p2_add_59901_comb;
  wire [31:0] p2_add_59894_comb;
  wire [31:0] p2_add_59895_comb;
  wire [31:0] p2_add_59896_comb;
  wire [31:0] p2_add_59897_comb;
  wire [31:0] p2_add_59890_comb;
  wire [31:0] p2_add_59891_comb;
  wire [31:0] p2_add_59892_comb;
  wire [31:0] p2_add_59893_comb;
  wire [31:0] p2_add_59886_comb;
  wire [31:0] p2_add_59887_comb;
  wire [31:0] p2_add_59888_comb;
  wire [31:0] p2_add_59889_comb;
  wire [31:0] p2_add_59882_comb;
  wire [31:0] p2_add_59883_comb;
  wire [31:0] p2_add_59884_comb;
  wire [31:0] p2_add_59885_comb;
  wire [31:0] p2_add_59878_comb;
  wire [31:0] p2_add_59879_comb;
  wire [31:0] p2_add_59880_comb;
  wire [31:0] p2_add_59881_comb;
  wire [31:0] p2_add_59874_comb;
  wire [31:0] p2_add_59875_comb;
  wire [31:0] p2_add_59876_comb;
  wire [31:0] p2_add_59877_comb;
  assign p2_smul_59866_comb = smul32b_32b_x_32b(p1_array_index_59094, p1_array_index_59038);
  assign p2_smul_59867_comb = smul32b_32b_x_32b(p1_array_index_59095, p1_array_index_59039);
  assign p2_smul_59868_comb = smul32b_32b_x_32b(p1_array_index_59096, p1_array_index_59040);
  assign p2_smul_59869_comb = smul32b_32b_x_32b(p1_array_index_59097, p1_array_index_59041);
  assign p2_smul_59870_comb = smul32b_32b_x_32b(p1_array_index_59098, p1_array_index_59042);
  assign p2_smul_59871_comb = smul32b_32b_x_32b(p1_array_index_59099, p1_array_index_59043);
  assign p2_smul_59872_comb = smul32b_32b_x_32b(p1_array_index_59100, p1_array_index_59044);
  assign p2_smul_59873_comb = smul32b_32b_x_32b(p1_array_index_59101, p1_array_index_59045);
  assign p2_smul_59858_comb = smul32b_32b_x_32b(p1_array_index_59094, p1_array_index_59030);
  assign p2_smul_59859_comb = smul32b_32b_x_32b(p1_array_index_59095, p1_array_index_59031);
  assign p2_smul_59860_comb = smul32b_32b_x_32b(p1_array_index_59096, p1_array_index_59032);
  assign p2_smul_59861_comb = smul32b_32b_x_32b(p1_array_index_59097, p1_array_index_59033);
  assign p2_smul_59862_comb = smul32b_32b_x_32b(p1_array_index_59098, p1_array_index_59034);
  assign p2_smul_59863_comb = smul32b_32b_x_32b(p1_array_index_59099, p1_array_index_59035);
  assign p2_smul_59864_comb = smul32b_32b_x_32b(p1_array_index_59100, p1_array_index_59036);
  assign p2_smul_59865_comb = smul32b_32b_x_32b(p1_array_index_59101, p1_array_index_59037);
  assign p2_smul_59850_comb = smul32b_32b_x_32b(p1_array_index_59094, p1_array_index_59022);
  assign p2_smul_59851_comb = smul32b_32b_x_32b(p1_array_index_59095, p1_array_index_59023);
  assign p2_smul_59852_comb = smul32b_32b_x_32b(p1_array_index_59096, p1_array_index_59024);
  assign p2_smul_59853_comb = smul32b_32b_x_32b(p1_array_index_59097, p1_array_index_59025);
  assign p2_smul_59854_comb = smul32b_32b_x_32b(p1_array_index_59098, p1_array_index_59026);
  assign p2_smul_59855_comb = smul32b_32b_x_32b(p1_array_index_59099, p1_array_index_59027);
  assign p2_smul_59856_comb = smul32b_32b_x_32b(p1_array_index_59100, p1_array_index_59028);
  assign p2_smul_59857_comb = smul32b_32b_x_32b(p1_array_index_59101, p1_array_index_59029);
  assign p2_smul_59842_comb = smul32b_32b_x_32b(p1_array_index_59094, p1_array_index_59014);
  assign p2_smul_59843_comb = smul32b_32b_x_32b(p1_array_index_59095, p1_array_index_59015);
  assign p2_smul_59844_comb = smul32b_32b_x_32b(p1_array_index_59096, p1_array_index_59016);
  assign p2_smul_59845_comb = smul32b_32b_x_32b(p1_array_index_59097, p1_array_index_59017);
  assign p2_smul_59846_comb = smul32b_32b_x_32b(p1_array_index_59098, p1_array_index_59018);
  assign p2_smul_59847_comb = smul32b_32b_x_32b(p1_array_index_59099, p1_array_index_59019);
  assign p2_smul_59848_comb = smul32b_32b_x_32b(p1_array_index_59100, p1_array_index_59020);
  assign p2_smul_59849_comb = smul32b_32b_x_32b(p1_array_index_59101, p1_array_index_59021);
  assign p2_smul_59834_comb = smul32b_32b_x_32b(p1_array_index_59094, p1_array_index_59006);
  assign p2_smul_59835_comb = smul32b_32b_x_32b(p1_array_index_59095, p1_array_index_59007);
  assign p2_smul_59836_comb = smul32b_32b_x_32b(p1_array_index_59096, p1_array_index_59008);
  assign p2_smul_59837_comb = smul32b_32b_x_32b(p1_array_index_59097, p1_array_index_59009);
  assign p2_smul_59838_comb = smul32b_32b_x_32b(p1_array_index_59098, p1_array_index_59010);
  assign p2_smul_59839_comb = smul32b_32b_x_32b(p1_array_index_59099, p1_array_index_59011);
  assign p2_smul_59840_comb = smul32b_32b_x_32b(p1_array_index_59100, p1_array_index_59012);
  assign p2_smul_59841_comb = smul32b_32b_x_32b(p1_array_index_59101, p1_array_index_59013);
  assign p2_smul_59826_comb = smul32b_32b_x_32b(p1_array_index_59094, p1_array_index_58998);
  assign p2_smul_59827_comb = smul32b_32b_x_32b(p1_array_index_59095, p1_array_index_58999);
  assign p2_smul_59828_comb = smul32b_32b_x_32b(p1_array_index_59096, p1_array_index_59000);
  assign p2_smul_59829_comb = smul32b_32b_x_32b(p1_array_index_59097, p1_array_index_59001);
  assign p2_smul_59830_comb = smul32b_32b_x_32b(p1_array_index_59098, p1_array_index_59002);
  assign p2_smul_59831_comb = smul32b_32b_x_32b(p1_array_index_59099, p1_array_index_59003);
  assign p2_smul_59832_comb = smul32b_32b_x_32b(p1_array_index_59100, p1_array_index_59004);
  assign p2_smul_59833_comb = smul32b_32b_x_32b(p1_array_index_59101, p1_array_index_59005);
  assign p2_smul_59818_comb = smul32b_32b_x_32b(p1_array_index_59094, p1_array_index_58990);
  assign p2_smul_59819_comb = smul32b_32b_x_32b(p1_array_index_59095, p1_array_index_58991);
  assign p2_smul_59820_comb = smul32b_32b_x_32b(p1_array_index_59096, p1_array_index_58992);
  assign p2_smul_59821_comb = smul32b_32b_x_32b(p1_array_index_59097, p1_array_index_58993);
  assign p2_smul_59822_comb = smul32b_32b_x_32b(p1_array_index_59098, p1_array_index_58994);
  assign p2_smul_59823_comb = smul32b_32b_x_32b(p1_array_index_59099, p1_array_index_58995);
  assign p2_smul_59824_comb = smul32b_32b_x_32b(p1_array_index_59100, p1_array_index_58996);
  assign p2_smul_59825_comb = smul32b_32b_x_32b(p1_array_index_59101, p1_array_index_58997);
  assign p2_smul_59810_comb = smul32b_32b_x_32b(p1_array_index_59094, p1_array_index_58975);
  assign p2_smul_59811_comb = smul32b_32b_x_32b(p1_array_index_59095, p1_array_index_58977);
  assign p2_smul_59812_comb = smul32b_32b_x_32b(p1_array_index_59096, p1_array_index_58979);
  assign p2_smul_59813_comb = smul32b_32b_x_32b(p1_array_index_59097, p1_array_index_58981);
  assign p2_smul_59814_comb = smul32b_32b_x_32b(p1_array_index_59098, p1_array_index_58983);
  assign p2_smul_59815_comb = smul32b_32b_x_32b(p1_array_index_59099, p1_array_index_58985);
  assign p2_smul_59816_comb = smul32b_32b_x_32b(p1_array_index_59100, p1_array_index_58987);
  assign p2_smul_59817_comb = smul32b_32b_x_32b(p1_array_index_59101, p1_array_index_58989);
  assign p2_smul_59802_comb = smul32b_32b_x_32b(p1_array_index_59086, p1_array_index_59038);
  assign p2_smul_59803_comb = smul32b_32b_x_32b(p1_array_index_59087, p1_array_index_59039);
  assign p2_smul_59804_comb = smul32b_32b_x_32b(p1_array_index_59088, p1_array_index_59040);
  assign p2_smul_59805_comb = smul32b_32b_x_32b(p1_array_index_59089, p1_array_index_59041);
  assign p2_smul_59806_comb = smul32b_32b_x_32b(p1_array_index_59090, p1_array_index_59042);
  assign p2_smul_59807_comb = smul32b_32b_x_32b(p1_array_index_59091, p1_array_index_59043);
  assign p2_smul_59808_comb = smul32b_32b_x_32b(p1_array_index_59092, p1_array_index_59044);
  assign p2_smul_59809_comb = smul32b_32b_x_32b(p1_array_index_59093, p1_array_index_59045);
  assign p2_smul_59794_comb = smul32b_32b_x_32b(p1_array_index_59086, p1_array_index_59030);
  assign p2_smul_59795_comb = smul32b_32b_x_32b(p1_array_index_59087, p1_array_index_59031);
  assign p2_smul_59796_comb = smul32b_32b_x_32b(p1_array_index_59088, p1_array_index_59032);
  assign p2_smul_59797_comb = smul32b_32b_x_32b(p1_array_index_59089, p1_array_index_59033);
  assign p2_smul_59798_comb = smul32b_32b_x_32b(p1_array_index_59090, p1_array_index_59034);
  assign p2_smul_59799_comb = smul32b_32b_x_32b(p1_array_index_59091, p1_array_index_59035);
  assign p2_smul_59800_comb = smul32b_32b_x_32b(p1_array_index_59092, p1_array_index_59036);
  assign p2_smul_59801_comb = smul32b_32b_x_32b(p1_array_index_59093, p1_array_index_59037);
  assign p2_smul_59786_comb = smul32b_32b_x_32b(p1_array_index_59086, p1_array_index_59022);
  assign p2_smul_59787_comb = smul32b_32b_x_32b(p1_array_index_59087, p1_array_index_59023);
  assign p2_smul_59788_comb = smul32b_32b_x_32b(p1_array_index_59088, p1_array_index_59024);
  assign p2_smul_59789_comb = smul32b_32b_x_32b(p1_array_index_59089, p1_array_index_59025);
  assign p2_smul_59790_comb = smul32b_32b_x_32b(p1_array_index_59090, p1_array_index_59026);
  assign p2_smul_59791_comb = smul32b_32b_x_32b(p1_array_index_59091, p1_array_index_59027);
  assign p2_smul_59792_comb = smul32b_32b_x_32b(p1_array_index_59092, p1_array_index_59028);
  assign p2_smul_59793_comb = smul32b_32b_x_32b(p1_array_index_59093, p1_array_index_59029);
  assign p2_smul_59778_comb = smul32b_32b_x_32b(p1_array_index_59086, p1_array_index_59014);
  assign p2_smul_59779_comb = smul32b_32b_x_32b(p1_array_index_59087, p1_array_index_59015);
  assign p2_smul_59780_comb = smul32b_32b_x_32b(p1_array_index_59088, p1_array_index_59016);
  assign p2_smul_59781_comb = smul32b_32b_x_32b(p1_array_index_59089, p1_array_index_59017);
  assign p2_smul_59782_comb = smul32b_32b_x_32b(p1_array_index_59090, p1_array_index_59018);
  assign p2_smul_59783_comb = smul32b_32b_x_32b(p1_array_index_59091, p1_array_index_59019);
  assign p2_smul_59784_comb = smul32b_32b_x_32b(p1_array_index_59092, p1_array_index_59020);
  assign p2_smul_59785_comb = smul32b_32b_x_32b(p1_array_index_59093, p1_array_index_59021);
  assign p2_smul_59770_comb = smul32b_32b_x_32b(p1_array_index_59086, p1_array_index_59006);
  assign p2_smul_59771_comb = smul32b_32b_x_32b(p1_array_index_59087, p1_array_index_59007);
  assign p2_smul_59772_comb = smul32b_32b_x_32b(p1_array_index_59088, p1_array_index_59008);
  assign p2_smul_59773_comb = smul32b_32b_x_32b(p1_array_index_59089, p1_array_index_59009);
  assign p2_smul_59774_comb = smul32b_32b_x_32b(p1_array_index_59090, p1_array_index_59010);
  assign p2_smul_59775_comb = smul32b_32b_x_32b(p1_array_index_59091, p1_array_index_59011);
  assign p2_smul_59776_comb = smul32b_32b_x_32b(p1_array_index_59092, p1_array_index_59012);
  assign p2_smul_59777_comb = smul32b_32b_x_32b(p1_array_index_59093, p1_array_index_59013);
  assign p2_smul_59762_comb = smul32b_32b_x_32b(p1_array_index_59086, p1_array_index_58998);
  assign p2_smul_59763_comb = smul32b_32b_x_32b(p1_array_index_59087, p1_array_index_58999);
  assign p2_smul_59764_comb = smul32b_32b_x_32b(p1_array_index_59088, p1_array_index_59000);
  assign p2_smul_59765_comb = smul32b_32b_x_32b(p1_array_index_59089, p1_array_index_59001);
  assign p2_smul_59766_comb = smul32b_32b_x_32b(p1_array_index_59090, p1_array_index_59002);
  assign p2_smul_59767_comb = smul32b_32b_x_32b(p1_array_index_59091, p1_array_index_59003);
  assign p2_smul_59768_comb = smul32b_32b_x_32b(p1_array_index_59092, p1_array_index_59004);
  assign p2_smul_59769_comb = smul32b_32b_x_32b(p1_array_index_59093, p1_array_index_59005);
  assign p2_smul_59754_comb = smul32b_32b_x_32b(p1_array_index_59086, p1_array_index_58990);
  assign p2_smul_59755_comb = smul32b_32b_x_32b(p1_array_index_59087, p1_array_index_58991);
  assign p2_smul_59756_comb = smul32b_32b_x_32b(p1_array_index_59088, p1_array_index_58992);
  assign p2_smul_59757_comb = smul32b_32b_x_32b(p1_array_index_59089, p1_array_index_58993);
  assign p2_smul_59758_comb = smul32b_32b_x_32b(p1_array_index_59090, p1_array_index_58994);
  assign p2_smul_59759_comb = smul32b_32b_x_32b(p1_array_index_59091, p1_array_index_58995);
  assign p2_smul_59760_comb = smul32b_32b_x_32b(p1_array_index_59092, p1_array_index_58996);
  assign p2_smul_59761_comb = smul32b_32b_x_32b(p1_array_index_59093, p1_array_index_58997);
  assign p2_smul_59746_comb = smul32b_32b_x_32b(p1_array_index_59086, p1_array_index_58975);
  assign p2_smul_59747_comb = smul32b_32b_x_32b(p1_array_index_59087, p1_array_index_58977);
  assign p2_smul_59748_comb = smul32b_32b_x_32b(p1_array_index_59088, p1_array_index_58979);
  assign p2_smul_59749_comb = smul32b_32b_x_32b(p1_array_index_59089, p1_array_index_58981);
  assign p2_smul_59750_comb = smul32b_32b_x_32b(p1_array_index_59090, p1_array_index_58983);
  assign p2_smul_59751_comb = smul32b_32b_x_32b(p1_array_index_59091, p1_array_index_58985);
  assign p2_smul_59752_comb = smul32b_32b_x_32b(p1_array_index_59092, p1_array_index_58987);
  assign p2_smul_59753_comb = smul32b_32b_x_32b(p1_array_index_59093, p1_array_index_58989);
  assign p2_smul_59738_comb = smul32b_32b_x_32b(p1_array_index_59078, p1_array_index_59038);
  assign p2_smul_59739_comb = smul32b_32b_x_32b(p1_array_index_59079, p1_array_index_59039);
  assign p2_smul_59740_comb = smul32b_32b_x_32b(p1_array_index_59080, p1_array_index_59040);
  assign p2_smul_59741_comb = smul32b_32b_x_32b(p1_array_index_59081, p1_array_index_59041);
  assign p2_smul_59742_comb = smul32b_32b_x_32b(p1_array_index_59082, p1_array_index_59042);
  assign p2_smul_59743_comb = smul32b_32b_x_32b(p1_array_index_59083, p1_array_index_59043);
  assign p2_smul_59744_comb = smul32b_32b_x_32b(p1_array_index_59084, p1_array_index_59044);
  assign p2_smul_59745_comb = smul32b_32b_x_32b(p1_array_index_59085, p1_array_index_59045);
  assign p2_smul_59730_comb = smul32b_32b_x_32b(p1_array_index_59078, p1_array_index_59030);
  assign p2_smul_59731_comb = smul32b_32b_x_32b(p1_array_index_59079, p1_array_index_59031);
  assign p2_smul_59732_comb = smul32b_32b_x_32b(p1_array_index_59080, p1_array_index_59032);
  assign p2_smul_59733_comb = smul32b_32b_x_32b(p1_array_index_59081, p1_array_index_59033);
  assign p2_smul_59734_comb = smul32b_32b_x_32b(p1_array_index_59082, p1_array_index_59034);
  assign p2_smul_59735_comb = smul32b_32b_x_32b(p1_array_index_59083, p1_array_index_59035);
  assign p2_smul_59736_comb = smul32b_32b_x_32b(p1_array_index_59084, p1_array_index_59036);
  assign p2_smul_59737_comb = smul32b_32b_x_32b(p1_array_index_59085, p1_array_index_59037);
  assign p2_smul_59722_comb = smul32b_32b_x_32b(p1_array_index_59078, p1_array_index_59022);
  assign p2_smul_59723_comb = smul32b_32b_x_32b(p1_array_index_59079, p1_array_index_59023);
  assign p2_smul_59724_comb = smul32b_32b_x_32b(p1_array_index_59080, p1_array_index_59024);
  assign p2_smul_59725_comb = smul32b_32b_x_32b(p1_array_index_59081, p1_array_index_59025);
  assign p2_smul_59726_comb = smul32b_32b_x_32b(p1_array_index_59082, p1_array_index_59026);
  assign p2_smul_59727_comb = smul32b_32b_x_32b(p1_array_index_59083, p1_array_index_59027);
  assign p2_smul_59728_comb = smul32b_32b_x_32b(p1_array_index_59084, p1_array_index_59028);
  assign p2_smul_59729_comb = smul32b_32b_x_32b(p1_array_index_59085, p1_array_index_59029);
  assign p2_smul_59714_comb = smul32b_32b_x_32b(p1_array_index_59078, p1_array_index_59014);
  assign p2_smul_59715_comb = smul32b_32b_x_32b(p1_array_index_59079, p1_array_index_59015);
  assign p2_smul_59716_comb = smul32b_32b_x_32b(p1_array_index_59080, p1_array_index_59016);
  assign p2_smul_59717_comb = smul32b_32b_x_32b(p1_array_index_59081, p1_array_index_59017);
  assign p2_smul_59718_comb = smul32b_32b_x_32b(p1_array_index_59082, p1_array_index_59018);
  assign p2_smul_59719_comb = smul32b_32b_x_32b(p1_array_index_59083, p1_array_index_59019);
  assign p2_smul_59720_comb = smul32b_32b_x_32b(p1_array_index_59084, p1_array_index_59020);
  assign p2_smul_59721_comb = smul32b_32b_x_32b(p1_array_index_59085, p1_array_index_59021);
  assign p2_smul_59706_comb = smul32b_32b_x_32b(p1_array_index_59078, p1_array_index_59006);
  assign p2_smul_59707_comb = smul32b_32b_x_32b(p1_array_index_59079, p1_array_index_59007);
  assign p2_smul_59708_comb = smul32b_32b_x_32b(p1_array_index_59080, p1_array_index_59008);
  assign p2_smul_59709_comb = smul32b_32b_x_32b(p1_array_index_59081, p1_array_index_59009);
  assign p2_smul_59710_comb = smul32b_32b_x_32b(p1_array_index_59082, p1_array_index_59010);
  assign p2_smul_59711_comb = smul32b_32b_x_32b(p1_array_index_59083, p1_array_index_59011);
  assign p2_smul_59712_comb = smul32b_32b_x_32b(p1_array_index_59084, p1_array_index_59012);
  assign p2_smul_59713_comb = smul32b_32b_x_32b(p1_array_index_59085, p1_array_index_59013);
  assign p2_smul_59698_comb = smul32b_32b_x_32b(p1_array_index_59078, p1_array_index_58998);
  assign p2_smul_59699_comb = smul32b_32b_x_32b(p1_array_index_59079, p1_array_index_58999);
  assign p2_smul_59700_comb = smul32b_32b_x_32b(p1_array_index_59080, p1_array_index_59000);
  assign p2_smul_59701_comb = smul32b_32b_x_32b(p1_array_index_59081, p1_array_index_59001);
  assign p2_smul_59702_comb = smul32b_32b_x_32b(p1_array_index_59082, p1_array_index_59002);
  assign p2_smul_59703_comb = smul32b_32b_x_32b(p1_array_index_59083, p1_array_index_59003);
  assign p2_smul_59704_comb = smul32b_32b_x_32b(p1_array_index_59084, p1_array_index_59004);
  assign p2_smul_59705_comb = smul32b_32b_x_32b(p1_array_index_59085, p1_array_index_59005);
  assign p2_smul_59690_comb = smul32b_32b_x_32b(p1_array_index_59078, p1_array_index_58990);
  assign p2_smul_59691_comb = smul32b_32b_x_32b(p1_array_index_59079, p1_array_index_58991);
  assign p2_smul_59692_comb = smul32b_32b_x_32b(p1_array_index_59080, p1_array_index_58992);
  assign p2_smul_59693_comb = smul32b_32b_x_32b(p1_array_index_59081, p1_array_index_58993);
  assign p2_smul_59694_comb = smul32b_32b_x_32b(p1_array_index_59082, p1_array_index_58994);
  assign p2_smul_59695_comb = smul32b_32b_x_32b(p1_array_index_59083, p1_array_index_58995);
  assign p2_smul_59696_comb = smul32b_32b_x_32b(p1_array_index_59084, p1_array_index_58996);
  assign p2_smul_59697_comb = smul32b_32b_x_32b(p1_array_index_59085, p1_array_index_58997);
  assign p2_smul_59682_comb = smul32b_32b_x_32b(p1_array_index_59078, p1_array_index_58975);
  assign p2_smul_59683_comb = smul32b_32b_x_32b(p1_array_index_59079, p1_array_index_58977);
  assign p2_smul_59684_comb = smul32b_32b_x_32b(p1_array_index_59080, p1_array_index_58979);
  assign p2_smul_59685_comb = smul32b_32b_x_32b(p1_array_index_59081, p1_array_index_58981);
  assign p2_smul_59686_comb = smul32b_32b_x_32b(p1_array_index_59082, p1_array_index_58983);
  assign p2_smul_59687_comb = smul32b_32b_x_32b(p1_array_index_59083, p1_array_index_58985);
  assign p2_smul_59688_comb = smul32b_32b_x_32b(p1_array_index_59084, p1_array_index_58987);
  assign p2_smul_59689_comb = smul32b_32b_x_32b(p1_array_index_59085, p1_array_index_58989);
  assign p2_smul_59674_comb = smul32b_32b_x_32b(p1_array_index_59070, p1_array_index_59038);
  assign p2_smul_59675_comb = smul32b_32b_x_32b(p1_array_index_59071, p1_array_index_59039);
  assign p2_smul_59676_comb = smul32b_32b_x_32b(p1_array_index_59072, p1_array_index_59040);
  assign p2_smul_59677_comb = smul32b_32b_x_32b(p1_array_index_59073, p1_array_index_59041);
  assign p2_smul_59678_comb = smul32b_32b_x_32b(p1_array_index_59074, p1_array_index_59042);
  assign p2_smul_59679_comb = smul32b_32b_x_32b(p1_array_index_59075, p1_array_index_59043);
  assign p2_smul_59680_comb = smul32b_32b_x_32b(p1_array_index_59076, p1_array_index_59044);
  assign p2_smul_59681_comb = smul32b_32b_x_32b(p1_array_index_59077, p1_array_index_59045);
  assign p2_smul_59666_comb = smul32b_32b_x_32b(p1_array_index_59070, p1_array_index_59030);
  assign p2_smul_59667_comb = smul32b_32b_x_32b(p1_array_index_59071, p1_array_index_59031);
  assign p2_smul_59668_comb = smul32b_32b_x_32b(p1_array_index_59072, p1_array_index_59032);
  assign p2_smul_59669_comb = smul32b_32b_x_32b(p1_array_index_59073, p1_array_index_59033);
  assign p2_smul_59670_comb = smul32b_32b_x_32b(p1_array_index_59074, p1_array_index_59034);
  assign p2_smul_59671_comb = smul32b_32b_x_32b(p1_array_index_59075, p1_array_index_59035);
  assign p2_smul_59672_comb = smul32b_32b_x_32b(p1_array_index_59076, p1_array_index_59036);
  assign p2_smul_59673_comb = smul32b_32b_x_32b(p1_array_index_59077, p1_array_index_59037);
  assign p2_smul_59658_comb = smul32b_32b_x_32b(p1_array_index_59070, p1_array_index_59022);
  assign p2_smul_59659_comb = smul32b_32b_x_32b(p1_array_index_59071, p1_array_index_59023);
  assign p2_smul_59660_comb = smul32b_32b_x_32b(p1_array_index_59072, p1_array_index_59024);
  assign p2_smul_59661_comb = smul32b_32b_x_32b(p1_array_index_59073, p1_array_index_59025);
  assign p2_smul_59662_comb = smul32b_32b_x_32b(p1_array_index_59074, p1_array_index_59026);
  assign p2_smul_59663_comb = smul32b_32b_x_32b(p1_array_index_59075, p1_array_index_59027);
  assign p2_smul_59664_comb = smul32b_32b_x_32b(p1_array_index_59076, p1_array_index_59028);
  assign p2_smul_59665_comb = smul32b_32b_x_32b(p1_array_index_59077, p1_array_index_59029);
  assign p2_smul_59650_comb = smul32b_32b_x_32b(p1_array_index_59070, p1_array_index_59014);
  assign p2_smul_59651_comb = smul32b_32b_x_32b(p1_array_index_59071, p1_array_index_59015);
  assign p2_smul_59652_comb = smul32b_32b_x_32b(p1_array_index_59072, p1_array_index_59016);
  assign p2_smul_59653_comb = smul32b_32b_x_32b(p1_array_index_59073, p1_array_index_59017);
  assign p2_smul_59654_comb = smul32b_32b_x_32b(p1_array_index_59074, p1_array_index_59018);
  assign p2_smul_59655_comb = smul32b_32b_x_32b(p1_array_index_59075, p1_array_index_59019);
  assign p2_smul_59656_comb = smul32b_32b_x_32b(p1_array_index_59076, p1_array_index_59020);
  assign p2_smul_59657_comb = smul32b_32b_x_32b(p1_array_index_59077, p1_array_index_59021);
  assign p2_smul_59642_comb = smul32b_32b_x_32b(p1_array_index_59070, p1_array_index_59006);
  assign p2_smul_59643_comb = smul32b_32b_x_32b(p1_array_index_59071, p1_array_index_59007);
  assign p2_smul_59644_comb = smul32b_32b_x_32b(p1_array_index_59072, p1_array_index_59008);
  assign p2_smul_59645_comb = smul32b_32b_x_32b(p1_array_index_59073, p1_array_index_59009);
  assign p2_smul_59646_comb = smul32b_32b_x_32b(p1_array_index_59074, p1_array_index_59010);
  assign p2_smul_59647_comb = smul32b_32b_x_32b(p1_array_index_59075, p1_array_index_59011);
  assign p2_smul_59648_comb = smul32b_32b_x_32b(p1_array_index_59076, p1_array_index_59012);
  assign p2_smul_59649_comb = smul32b_32b_x_32b(p1_array_index_59077, p1_array_index_59013);
  assign p2_smul_59634_comb = smul32b_32b_x_32b(p1_array_index_59070, p1_array_index_58998);
  assign p2_smul_59635_comb = smul32b_32b_x_32b(p1_array_index_59071, p1_array_index_58999);
  assign p2_smul_59636_comb = smul32b_32b_x_32b(p1_array_index_59072, p1_array_index_59000);
  assign p2_smul_59637_comb = smul32b_32b_x_32b(p1_array_index_59073, p1_array_index_59001);
  assign p2_smul_59638_comb = smul32b_32b_x_32b(p1_array_index_59074, p1_array_index_59002);
  assign p2_smul_59639_comb = smul32b_32b_x_32b(p1_array_index_59075, p1_array_index_59003);
  assign p2_smul_59640_comb = smul32b_32b_x_32b(p1_array_index_59076, p1_array_index_59004);
  assign p2_smul_59641_comb = smul32b_32b_x_32b(p1_array_index_59077, p1_array_index_59005);
  assign p2_smul_59626_comb = smul32b_32b_x_32b(p1_array_index_59070, p1_array_index_58990);
  assign p2_smul_59627_comb = smul32b_32b_x_32b(p1_array_index_59071, p1_array_index_58991);
  assign p2_smul_59628_comb = smul32b_32b_x_32b(p1_array_index_59072, p1_array_index_58992);
  assign p2_smul_59629_comb = smul32b_32b_x_32b(p1_array_index_59073, p1_array_index_58993);
  assign p2_smul_59630_comb = smul32b_32b_x_32b(p1_array_index_59074, p1_array_index_58994);
  assign p2_smul_59631_comb = smul32b_32b_x_32b(p1_array_index_59075, p1_array_index_58995);
  assign p2_smul_59632_comb = smul32b_32b_x_32b(p1_array_index_59076, p1_array_index_58996);
  assign p2_smul_59633_comb = smul32b_32b_x_32b(p1_array_index_59077, p1_array_index_58997);
  assign p2_smul_59618_comb = smul32b_32b_x_32b(p1_array_index_59070, p1_array_index_58975);
  assign p2_smul_59619_comb = smul32b_32b_x_32b(p1_array_index_59071, p1_array_index_58977);
  assign p2_smul_59620_comb = smul32b_32b_x_32b(p1_array_index_59072, p1_array_index_58979);
  assign p2_smul_59621_comb = smul32b_32b_x_32b(p1_array_index_59073, p1_array_index_58981);
  assign p2_smul_59622_comb = smul32b_32b_x_32b(p1_array_index_59074, p1_array_index_58983);
  assign p2_smul_59623_comb = smul32b_32b_x_32b(p1_array_index_59075, p1_array_index_58985);
  assign p2_smul_59624_comb = smul32b_32b_x_32b(p1_array_index_59076, p1_array_index_58987);
  assign p2_smul_59625_comb = smul32b_32b_x_32b(p1_array_index_59077, p1_array_index_58989);
  assign p2_smul_59610_comb = smul32b_32b_x_32b(p1_array_index_59062, p1_array_index_59038);
  assign p2_smul_59611_comb = smul32b_32b_x_32b(p1_array_index_59063, p1_array_index_59039);
  assign p2_smul_59612_comb = smul32b_32b_x_32b(p1_array_index_59064, p1_array_index_59040);
  assign p2_smul_59613_comb = smul32b_32b_x_32b(p1_array_index_59065, p1_array_index_59041);
  assign p2_smul_59614_comb = smul32b_32b_x_32b(p1_array_index_59066, p1_array_index_59042);
  assign p2_smul_59615_comb = smul32b_32b_x_32b(p1_array_index_59067, p1_array_index_59043);
  assign p2_smul_59616_comb = smul32b_32b_x_32b(p1_array_index_59068, p1_array_index_59044);
  assign p2_smul_59617_comb = smul32b_32b_x_32b(p1_array_index_59069, p1_array_index_59045);
  assign p2_smul_59602_comb = smul32b_32b_x_32b(p1_array_index_59062, p1_array_index_59030);
  assign p2_smul_59603_comb = smul32b_32b_x_32b(p1_array_index_59063, p1_array_index_59031);
  assign p2_smul_59604_comb = smul32b_32b_x_32b(p1_array_index_59064, p1_array_index_59032);
  assign p2_smul_59605_comb = smul32b_32b_x_32b(p1_array_index_59065, p1_array_index_59033);
  assign p2_smul_59606_comb = smul32b_32b_x_32b(p1_array_index_59066, p1_array_index_59034);
  assign p2_smul_59607_comb = smul32b_32b_x_32b(p1_array_index_59067, p1_array_index_59035);
  assign p2_smul_59608_comb = smul32b_32b_x_32b(p1_array_index_59068, p1_array_index_59036);
  assign p2_smul_59609_comb = smul32b_32b_x_32b(p1_array_index_59069, p1_array_index_59037);
  assign p2_smul_59594_comb = smul32b_32b_x_32b(p1_array_index_59062, p1_array_index_59022);
  assign p2_smul_59595_comb = smul32b_32b_x_32b(p1_array_index_59063, p1_array_index_59023);
  assign p2_smul_59596_comb = smul32b_32b_x_32b(p1_array_index_59064, p1_array_index_59024);
  assign p2_smul_59597_comb = smul32b_32b_x_32b(p1_array_index_59065, p1_array_index_59025);
  assign p2_smul_59598_comb = smul32b_32b_x_32b(p1_array_index_59066, p1_array_index_59026);
  assign p2_smul_59599_comb = smul32b_32b_x_32b(p1_array_index_59067, p1_array_index_59027);
  assign p2_smul_59600_comb = smul32b_32b_x_32b(p1_array_index_59068, p1_array_index_59028);
  assign p2_smul_59601_comb = smul32b_32b_x_32b(p1_array_index_59069, p1_array_index_59029);
  assign p2_smul_59586_comb = smul32b_32b_x_32b(p1_array_index_59062, p1_array_index_59014);
  assign p2_smul_59587_comb = smul32b_32b_x_32b(p1_array_index_59063, p1_array_index_59015);
  assign p2_smul_59588_comb = smul32b_32b_x_32b(p1_array_index_59064, p1_array_index_59016);
  assign p2_smul_59589_comb = smul32b_32b_x_32b(p1_array_index_59065, p1_array_index_59017);
  assign p2_smul_59590_comb = smul32b_32b_x_32b(p1_array_index_59066, p1_array_index_59018);
  assign p2_smul_59591_comb = smul32b_32b_x_32b(p1_array_index_59067, p1_array_index_59019);
  assign p2_smul_59592_comb = smul32b_32b_x_32b(p1_array_index_59068, p1_array_index_59020);
  assign p2_smul_59593_comb = smul32b_32b_x_32b(p1_array_index_59069, p1_array_index_59021);
  assign p2_smul_59578_comb = smul32b_32b_x_32b(p1_array_index_59062, p1_array_index_59006);
  assign p2_smul_59579_comb = smul32b_32b_x_32b(p1_array_index_59063, p1_array_index_59007);
  assign p2_smul_59580_comb = smul32b_32b_x_32b(p1_array_index_59064, p1_array_index_59008);
  assign p2_smul_59581_comb = smul32b_32b_x_32b(p1_array_index_59065, p1_array_index_59009);
  assign p2_smul_59582_comb = smul32b_32b_x_32b(p1_array_index_59066, p1_array_index_59010);
  assign p2_smul_59583_comb = smul32b_32b_x_32b(p1_array_index_59067, p1_array_index_59011);
  assign p2_smul_59584_comb = smul32b_32b_x_32b(p1_array_index_59068, p1_array_index_59012);
  assign p2_smul_59585_comb = smul32b_32b_x_32b(p1_array_index_59069, p1_array_index_59013);
  assign p2_smul_59570_comb = smul32b_32b_x_32b(p1_array_index_59062, p1_array_index_58998);
  assign p2_smul_59571_comb = smul32b_32b_x_32b(p1_array_index_59063, p1_array_index_58999);
  assign p2_smul_59572_comb = smul32b_32b_x_32b(p1_array_index_59064, p1_array_index_59000);
  assign p2_smul_59573_comb = smul32b_32b_x_32b(p1_array_index_59065, p1_array_index_59001);
  assign p2_smul_59574_comb = smul32b_32b_x_32b(p1_array_index_59066, p1_array_index_59002);
  assign p2_smul_59575_comb = smul32b_32b_x_32b(p1_array_index_59067, p1_array_index_59003);
  assign p2_smul_59576_comb = smul32b_32b_x_32b(p1_array_index_59068, p1_array_index_59004);
  assign p2_smul_59577_comb = smul32b_32b_x_32b(p1_array_index_59069, p1_array_index_59005);
  assign p2_smul_59562_comb = smul32b_32b_x_32b(p1_array_index_59062, p1_array_index_58990);
  assign p2_smul_59563_comb = smul32b_32b_x_32b(p1_array_index_59063, p1_array_index_58991);
  assign p2_smul_59564_comb = smul32b_32b_x_32b(p1_array_index_59064, p1_array_index_58992);
  assign p2_smul_59565_comb = smul32b_32b_x_32b(p1_array_index_59065, p1_array_index_58993);
  assign p2_smul_59566_comb = smul32b_32b_x_32b(p1_array_index_59066, p1_array_index_58994);
  assign p2_smul_59567_comb = smul32b_32b_x_32b(p1_array_index_59067, p1_array_index_58995);
  assign p2_smul_59568_comb = smul32b_32b_x_32b(p1_array_index_59068, p1_array_index_58996);
  assign p2_smul_59569_comb = smul32b_32b_x_32b(p1_array_index_59069, p1_array_index_58997);
  assign p2_smul_59554_comb = smul32b_32b_x_32b(p1_array_index_59062, p1_array_index_58975);
  assign p2_smul_59555_comb = smul32b_32b_x_32b(p1_array_index_59063, p1_array_index_58977);
  assign p2_smul_59556_comb = smul32b_32b_x_32b(p1_array_index_59064, p1_array_index_58979);
  assign p2_smul_59557_comb = smul32b_32b_x_32b(p1_array_index_59065, p1_array_index_58981);
  assign p2_smul_59558_comb = smul32b_32b_x_32b(p1_array_index_59066, p1_array_index_58983);
  assign p2_smul_59559_comb = smul32b_32b_x_32b(p1_array_index_59067, p1_array_index_58985);
  assign p2_smul_59560_comb = smul32b_32b_x_32b(p1_array_index_59068, p1_array_index_58987);
  assign p2_smul_59561_comb = smul32b_32b_x_32b(p1_array_index_59069, p1_array_index_58989);
  assign p2_smul_59546_comb = smul32b_32b_x_32b(p1_array_index_59054, p1_array_index_59038);
  assign p2_smul_59547_comb = smul32b_32b_x_32b(p1_array_index_59055, p1_array_index_59039);
  assign p2_smul_59548_comb = smul32b_32b_x_32b(p1_array_index_59056, p1_array_index_59040);
  assign p2_smul_59549_comb = smul32b_32b_x_32b(p1_array_index_59057, p1_array_index_59041);
  assign p2_smul_59550_comb = smul32b_32b_x_32b(p1_array_index_59058, p1_array_index_59042);
  assign p2_smul_59551_comb = smul32b_32b_x_32b(p1_array_index_59059, p1_array_index_59043);
  assign p2_smul_59552_comb = smul32b_32b_x_32b(p1_array_index_59060, p1_array_index_59044);
  assign p2_smul_59553_comb = smul32b_32b_x_32b(p1_array_index_59061, p1_array_index_59045);
  assign p2_smul_59538_comb = smul32b_32b_x_32b(p1_array_index_59054, p1_array_index_59030);
  assign p2_smul_59539_comb = smul32b_32b_x_32b(p1_array_index_59055, p1_array_index_59031);
  assign p2_smul_59540_comb = smul32b_32b_x_32b(p1_array_index_59056, p1_array_index_59032);
  assign p2_smul_59541_comb = smul32b_32b_x_32b(p1_array_index_59057, p1_array_index_59033);
  assign p2_smul_59542_comb = smul32b_32b_x_32b(p1_array_index_59058, p1_array_index_59034);
  assign p2_smul_59543_comb = smul32b_32b_x_32b(p1_array_index_59059, p1_array_index_59035);
  assign p2_smul_59544_comb = smul32b_32b_x_32b(p1_array_index_59060, p1_array_index_59036);
  assign p2_smul_59545_comb = smul32b_32b_x_32b(p1_array_index_59061, p1_array_index_59037);
  assign p2_smul_59530_comb = smul32b_32b_x_32b(p1_array_index_59054, p1_array_index_59022);
  assign p2_smul_59531_comb = smul32b_32b_x_32b(p1_array_index_59055, p1_array_index_59023);
  assign p2_smul_59532_comb = smul32b_32b_x_32b(p1_array_index_59056, p1_array_index_59024);
  assign p2_smul_59533_comb = smul32b_32b_x_32b(p1_array_index_59057, p1_array_index_59025);
  assign p2_smul_59534_comb = smul32b_32b_x_32b(p1_array_index_59058, p1_array_index_59026);
  assign p2_smul_59535_comb = smul32b_32b_x_32b(p1_array_index_59059, p1_array_index_59027);
  assign p2_smul_59536_comb = smul32b_32b_x_32b(p1_array_index_59060, p1_array_index_59028);
  assign p2_smul_59537_comb = smul32b_32b_x_32b(p1_array_index_59061, p1_array_index_59029);
  assign p2_smul_59522_comb = smul32b_32b_x_32b(p1_array_index_59054, p1_array_index_59014);
  assign p2_smul_59523_comb = smul32b_32b_x_32b(p1_array_index_59055, p1_array_index_59015);
  assign p2_smul_59524_comb = smul32b_32b_x_32b(p1_array_index_59056, p1_array_index_59016);
  assign p2_smul_59525_comb = smul32b_32b_x_32b(p1_array_index_59057, p1_array_index_59017);
  assign p2_smul_59526_comb = smul32b_32b_x_32b(p1_array_index_59058, p1_array_index_59018);
  assign p2_smul_59527_comb = smul32b_32b_x_32b(p1_array_index_59059, p1_array_index_59019);
  assign p2_smul_59528_comb = smul32b_32b_x_32b(p1_array_index_59060, p1_array_index_59020);
  assign p2_smul_59529_comb = smul32b_32b_x_32b(p1_array_index_59061, p1_array_index_59021);
  assign p2_smul_59514_comb = smul32b_32b_x_32b(p1_array_index_59054, p1_array_index_59006);
  assign p2_smul_59515_comb = smul32b_32b_x_32b(p1_array_index_59055, p1_array_index_59007);
  assign p2_smul_59516_comb = smul32b_32b_x_32b(p1_array_index_59056, p1_array_index_59008);
  assign p2_smul_59517_comb = smul32b_32b_x_32b(p1_array_index_59057, p1_array_index_59009);
  assign p2_smul_59518_comb = smul32b_32b_x_32b(p1_array_index_59058, p1_array_index_59010);
  assign p2_smul_59519_comb = smul32b_32b_x_32b(p1_array_index_59059, p1_array_index_59011);
  assign p2_smul_59520_comb = smul32b_32b_x_32b(p1_array_index_59060, p1_array_index_59012);
  assign p2_smul_59521_comb = smul32b_32b_x_32b(p1_array_index_59061, p1_array_index_59013);
  assign p2_smul_59506_comb = smul32b_32b_x_32b(p1_array_index_59054, p1_array_index_58998);
  assign p2_smul_59507_comb = smul32b_32b_x_32b(p1_array_index_59055, p1_array_index_58999);
  assign p2_smul_59508_comb = smul32b_32b_x_32b(p1_array_index_59056, p1_array_index_59000);
  assign p2_smul_59509_comb = smul32b_32b_x_32b(p1_array_index_59057, p1_array_index_59001);
  assign p2_smul_59510_comb = smul32b_32b_x_32b(p1_array_index_59058, p1_array_index_59002);
  assign p2_smul_59511_comb = smul32b_32b_x_32b(p1_array_index_59059, p1_array_index_59003);
  assign p2_smul_59512_comb = smul32b_32b_x_32b(p1_array_index_59060, p1_array_index_59004);
  assign p2_smul_59513_comb = smul32b_32b_x_32b(p1_array_index_59061, p1_array_index_59005);
  assign p2_smul_59498_comb = smul32b_32b_x_32b(p1_array_index_59054, p1_array_index_58990);
  assign p2_smul_59499_comb = smul32b_32b_x_32b(p1_array_index_59055, p1_array_index_58991);
  assign p2_smul_59500_comb = smul32b_32b_x_32b(p1_array_index_59056, p1_array_index_58992);
  assign p2_smul_59501_comb = smul32b_32b_x_32b(p1_array_index_59057, p1_array_index_58993);
  assign p2_smul_59502_comb = smul32b_32b_x_32b(p1_array_index_59058, p1_array_index_58994);
  assign p2_smul_59503_comb = smul32b_32b_x_32b(p1_array_index_59059, p1_array_index_58995);
  assign p2_smul_59504_comb = smul32b_32b_x_32b(p1_array_index_59060, p1_array_index_58996);
  assign p2_smul_59505_comb = smul32b_32b_x_32b(p1_array_index_59061, p1_array_index_58997);
  assign p2_smul_59490_comb = smul32b_32b_x_32b(p1_array_index_59054, p1_array_index_58975);
  assign p2_smul_59491_comb = smul32b_32b_x_32b(p1_array_index_59055, p1_array_index_58977);
  assign p2_smul_59492_comb = smul32b_32b_x_32b(p1_array_index_59056, p1_array_index_58979);
  assign p2_smul_59493_comb = smul32b_32b_x_32b(p1_array_index_59057, p1_array_index_58981);
  assign p2_smul_59494_comb = smul32b_32b_x_32b(p1_array_index_59058, p1_array_index_58983);
  assign p2_smul_59495_comb = smul32b_32b_x_32b(p1_array_index_59059, p1_array_index_58985);
  assign p2_smul_59496_comb = smul32b_32b_x_32b(p1_array_index_59060, p1_array_index_58987);
  assign p2_smul_59497_comb = smul32b_32b_x_32b(p1_array_index_59061, p1_array_index_58989);
  assign p2_smul_59482_comb = smul32b_32b_x_32b(p1_array_index_59046, p1_array_index_59038);
  assign p2_smul_59483_comb = smul32b_32b_x_32b(p1_array_index_59047, p1_array_index_59039);
  assign p2_smul_59484_comb = smul32b_32b_x_32b(p1_array_index_59048, p1_array_index_59040);
  assign p2_smul_59485_comb = smul32b_32b_x_32b(p1_array_index_59049, p1_array_index_59041);
  assign p2_smul_59486_comb = smul32b_32b_x_32b(p1_array_index_59050, p1_array_index_59042);
  assign p2_smul_59487_comb = smul32b_32b_x_32b(p1_array_index_59051, p1_array_index_59043);
  assign p2_smul_59488_comb = smul32b_32b_x_32b(p1_array_index_59052, p1_array_index_59044);
  assign p2_smul_59489_comb = smul32b_32b_x_32b(p1_array_index_59053, p1_array_index_59045);
  assign p2_smul_59474_comb = smul32b_32b_x_32b(p1_array_index_59046, p1_array_index_59030);
  assign p2_smul_59475_comb = smul32b_32b_x_32b(p1_array_index_59047, p1_array_index_59031);
  assign p2_smul_59476_comb = smul32b_32b_x_32b(p1_array_index_59048, p1_array_index_59032);
  assign p2_smul_59477_comb = smul32b_32b_x_32b(p1_array_index_59049, p1_array_index_59033);
  assign p2_smul_59478_comb = smul32b_32b_x_32b(p1_array_index_59050, p1_array_index_59034);
  assign p2_smul_59479_comb = smul32b_32b_x_32b(p1_array_index_59051, p1_array_index_59035);
  assign p2_smul_59480_comb = smul32b_32b_x_32b(p1_array_index_59052, p1_array_index_59036);
  assign p2_smul_59481_comb = smul32b_32b_x_32b(p1_array_index_59053, p1_array_index_59037);
  assign p2_smul_59466_comb = smul32b_32b_x_32b(p1_array_index_59046, p1_array_index_59022);
  assign p2_smul_59467_comb = smul32b_32b_x_32b(p1_array_index_59047, p1_array_index_59023);
  assign p2_smul_59468_comb = smul32b_32b_x_32b(p1_array_index_59048, p1_array_index_59024);
  assign p2_smul_59469_comb = smul32b_32b_x_32b(p1_array_index_59049, p1_array_index_59025);
  assign p2_smul_59470_comb = smul32b_32b_x_32b(p1_array_index_59050, p1_array_index_59026);
  assign p2_smul_59471_comb = smul32b_32b_x_32b(p1_array_index_59051, p1_array_index_59027);
  assign p2_smul_59472_comb = smul32b_32b_x_32b(p1_array_index_59052, p1_array_index_59028);
  assign p2_smul_59473_comb = smul32b_32b_x_32b(p1_array_index_59053, p1_array_index_59029);
  assign p2_smul_59458_comb = smul32b_32b_x_32b(p1_array_index_59046, p1_array_index_59014);
  assign p2_smul_59459_comb = smul32b_32b_x_32b(p1_array_index_59047, p1_array_index_59015);
  assign p2_smul_59460_comb = smul32b_32b_x_32b(p1_array_index_59048, p1_array_index_59016);
  assign p2_smul_59461_comb = smul32b_32b_x_32b(p1_array_index_59049, p1_array_index_59017);
  assign p2_smul_59462_comb = smul32b_32b_x_32b(p1_array_index_59050, p1_array_index_59018);
  assign p2_smul_59463_comb = smul32b_32b_x_32b(p1_array_index_59051, p1_array_index_59019);
  assign p2_smul_59464_comb = smul32b_32b_x_32b(p1_array_index_59052, p1_array_index_59020);
  assign p2_smul_59465_comb = smul32b_32b_x_32b(p1_array_index_59053, p1_array_index_59021);
  assign p2_smul_59450_comb = smul32b_32b_x_32b(p1_array_index_59046, p1_array_index_59006);
  assign p2_smul_59451_comb = smul32b_32b_x_32b(p1_array_index_59047, p1_array_index_59007);
  assign p2_smul_59452_comb = smul32b_32b_x_32b(p1_array_index_59048, p1_array_index_59008);
  assign p2_smul_59453_comb = smul32b_32b_x_32b(p1_array_index_59049, p1_array_index_59009);
  assign p2_smul_59454_comb = smul32b_32b_x_32b(p1_array_index_59050, p1_array_index_59010);
  assign p2_smul_59455_comb = smul32b_32b_x_32b(p1_array_index_59051, p1_array_index_59011);
  assign p2_smul_59456_comb = smul32b_32b_x_32b(p1_array_index_59052, p1_array_index_59012);
  assign p2_smul_59457_comb = smul32b_32b_x_32b(p1_array_index_59053, p1_array_index_59013);
  assign p2_smul_59442_comb = smul32b_32b_x_32b(p1_array_index_59046, p1_array_index_58998);
  assign p2_smul_59443_comb = smul32b_32b_x_32b(p1_array_index_59047, p1_array_index_58999);
  assign p2_smul_59444_comb = smul32b_32b_x_32b(p1_array_index_59048, p1_array_index_59000);
  assign p2_smul_59445_comb = smul32b_32b_x_32b(p1_array_index_59049, p1_array_index_59001);
  assign p2_smul_59446_comb = smul32b_32b_x_32b(p1_array_index_59050, p1_array_index_59002);
  assign p2_smul_59447_comb = smul32b_32b_x_32b(p1_array_index_59051, p1_array_index_59003);
  assign p2_smul_59448_comb = smul32b_32b_x_32b(p1_array_index_59052, p1_array_index_59004);
  assign p2_smul_59449_comb = smul32b_32b_x_32b(p1_array_index_59053, p1_array_index_59005);
  assign p2_smul_59434_comb = smul32b_32b_x_32b(p1_array_index_59046, p1_array_index_58990);
  assign p2_smul_59435_comb = smul32b_32b_x_32b(p1_array_index_59047, p1_array_index_58991);
  assign p2_smul_59436_comb = smul32b_32b_x_32b(p1_array_index_59048, p1_array_index_58992);
  assign p2_smul_59437_comb = smul32b_32b_x_32b(p1_array_index_59049, p1_array_index_58993);
  assign p2_smul_59438_comb = smul32b_32b_x_32b(p1_array_index_59050, p1_array_index_58994);
  assign p2_smul_59439_comb = smul32b_32b_x_32b(p1_array_index_59051, p1_array_index_58995);
  assign p2_smul_59440_comb = smul32b_32b_x_32b(p1_array_index_59052, p1_array_index_58996);
  assign p2_smul_59441_comb = smul32b_32b_x_32b(p1_array_index_59053, p1_array_index_58997);
  assign p2_smul_59426_comb = smul32b_32b_x_32b(p1_array_index_59046, p1_array_index_58975);
  assign p2_smul_59427_comb = smul32b_32b_x_32b(p1_array_index_59047, p1_array_index_58977);
  assign p2_smul_59428_comb = smul32b_32b_x_32b(p1_array_index_59048, p1_array_index_58979);
  assign p2_smul_59429_comb = smul32b_32b_x_32b(p1_array_index_59049, p1_array_index_58981);
  assign p2_smul_59430_comb = smul32b_32b_x_32b(p1_array_index_59050, p1_array_index_58983);
  assign p2_smul_59431_comb = smul32b_32b_x_32b(p1_array_index_59051, p1_array_index_58985);
  assign p2_smul_59432_comb = smul32b_32b_x_32b(p1_array_index_59052, p1_array_index_58987);
  assign p2_smul_59433_comb = smul32b_32b_x_32b(p1_array_index_59053, p1_array_index_58989);
  assign p2_smul_59418_comb = smul32b_32b_x_32b(p1_array_index_58974, p1_array_index_59038);
  assign p2_smul_59419_comb = smul32b_32b_x_32b(p1_array_index_58976, p1_array_index_59039);
  assign p2_smul_59420_comb = smul32b_32b_x_32b(p1_array_index_58978, p1_array_index_59040);
  assign p2_smul_59421_comb = smul32b_32b_x_32b(p1_array_index_58980, p1_array_index_59041);
  assign p2_smul_59422_comb = smul32b_32b_x_32b(p1_array_index_58982, p1_array_index_59042);
  assign p2_smul_59423_comb = smul32b_32b_x_32b(p1_array_index_58984, p1_array_index_59043);
  assign p2_smul_59424_comb = smul32b_32b_x_32b(p1_array_index_58986, p1_array_index_59044);
  assign p2_smul_59425_comb = smul32b_32b_x_32b(p1_array_index_58988, p1_array_index_59045);
  assign p2_smul_59410_comb = smul32b_32b_x_32b(p1_array_index_58974, p1_array_index_59030);
  assign p2_smul_59411_comb = smul32b_32b_x_32b(p1_array_index_58976, p1_array_index_59031);
  assign p2_smul_59412_comb = smul32b_32b_x_32b(p1_array_index_58978, p1_array_index_59032);
  assign p2_smul_59413_comb = smul32b_32b_x_32b(p1_array_index_58980, p1_array_index_59033);
  assign p2_smul_59414_comb = smul32b_32b_x_32b(p1_array_index_58982, p1_array_index_59034);
  assign p2_smul_59415_comb = smul32b_32b_x_32b(p1_array_index_58984, p1_array_index_59035);
  assign p2_smul_59416_comb = smul32b_32b_x_32b(p1_array_index_58986, p1_array_index_59036);
  assign p2_smul_59417_comb = smul32b_32b_x_32b(p1_array_index_58988, p1_array_index_59037);
  assign p2_smul_59402_comb = smul32b_32b_x_32b(p1_array_index_58974, p1_array_index_59022);
  assign p2_smul_59403_comb = smul32b_32b_x_32b(p1_array_index_58976, p1_array_index_59023);
  assign p2_smul_59404_comb = smul32b_32b_x_32b(p1_array_index_58978, p1_array_index_59024);
  assign p2_smul_59405_comb = smul32b_32b_x_32b(p1_array_index_58980, p1_array_index_59025);
  assign p2_smul_59406_comb = smul32b_32b_x_32b(p1_array_index_58982, p1_array_index_59026);
  assign p2_smul_59407_comb = smul32b_32b_x_32b(p1_array_index_58984, p1_array_index_59027);
  assign p2_smul_59408_comb = smul32b_32b_x_32b(p1_array_index_58986, p1_array_index_59028);
  assign p2_smul_59409_comb = smul32b_32b_x_32b(p1_array_index_58988, p1_array_index_59029);
  assign p2_smul_59394_comb = smul32b_32b_x_32b(p1_array_index_58974, p1_array_index_59014);
  assign p2_smul_59395_comb = smul32b_32b_x_32b(p1_array_index_58976, p1_array_index_59015);
  assign p2_smul_59396_comb = smul32b_32b_x_32b(p1_array_index_58978, p1_array_index_59016);
  assign p2_smul_59397_comb = smul32b_32b_x_32b(p1_array_index_58980, p1_array_index_59017);
  assign p2_smul_59398_comb = smul32b_32b_x_32b(p1_array_index_58982, p1_array_index_59018);
  assign p2_smul_59399_comb = smul32b_32b_x_32b(p1_array_index_58984, p1_array_index_59019);
  assign p2_smul_59400_comb = smul32b_32b_x_32b(p1_array_index_58986, p1_array_index_59020);
  assign p2_smul_59401_comb = smul32b_32b_x_32b(p1_array_index_58988, p1_array_index_59021);
  assign p2_smul_59386_comb = smul32b_32b_x_32b(p1_array_index_58974, p1_array_index_59006);
  assign p2_smul_59387_comb = smul32b_32b_x_32b(p1_array_index_58976, p1_array_index_59007);
  assign p2_smul_59388_comb = smul32b_32b_x_32b(p1_array_index_58978, p1_array_index_59008);
  assign p2_smul_59389_comb = smul32b_32b_x_32b(p1_array_index_58980, p1_array_index_59009);
  assign p2_smul_59390_comb = smul32b_32b_x_32b(p1_array_index_58982, p1_array_index_59010);
  assign p2_smul_59391_comb = smul32b_32b_x_32b(p1_array_index_58984, p1_array_index_59011);
  assign p2_smul_59392_comb = smul32b_32b_x_32b(p1_array_index_58986, p1_array_index_59012);
  assign p2_smul_59393_comb = smul32b_32b_x_32b(p1_array_index_58988, p1_array_index_59013);
  assign p2_smul_59378_comb = smul32b_32b_x_32b(p1_array_index_58974, p1_array_index_58998);
  assign p2_smul_59379_comb = smul32b_32b_x_32b(p1_array_index_58976, p1_array_index_58999);
  assign p2_smul_59380_comb = smul32b_32b_x_32b(p1_array_index_58978, p1_array_index_59000);
  assign p2_smul_59381_comb = smul32b_32b_x_32b(p1_array_index_58980, p1_array_index_59001);
  assign p2_smul_59382_comb = smul32b_32b_x_32b(p1_array_index_58982, p1_array_index_59002);
  assign p2_smul_59383_comb = smul32b_32b_x_32b(p1_array_index_58984, p1_array_index_59003);
  assign p2_smul_59384_comb = smul32b_32b_x_32b(p1_array_index_58986, p1_array_index_59004);
  assign p2_smul_59385_comb = smul32b_32b_x_32b(p1_array_index_58988, p1_array_index_59005);
  assign p2_smul_59370_comb = smul32b_32b_x_32b(p1_array_index_58974, p1_array_index_58990);
  assign p2_smul_59371_comb = smul32b_32b_x_32b(p1_array_index_58976, p1_array_index_58991);
  assign p2_smul_59372_comb = smul32b_32b_x_32b(p1_array_index_58978, p1_array_index_58992);
  assign p2_smul_59373_comb = smul32b_32b_x_32b(p1_array_index_58980, p1_array_index_58993);
  assign p2_smul_59374_comb = smul32b_32b_x_32b(p1_array_index_58982, p1_array_index_58994);
  assign p2_smul_59375_comb = smul32b_32b_x_32b(p1_array_index_58984, p1_array_index_58995);
  assign p2_smul_59376_comb = smul32b_32b_x_32b(p1_array_index_58986, p1_array_index_58996);
  assign p2_smul_59377_comb = smul32b_32b_x_32b(p1_array_index_58988, p1_array_index_58997);
  assign p2_smul_59362_comb = smul32b_32b_x_32b(p1_array_index_58974, p1_array_index_58975);
  assign p2_smul_59363_comb = smul32b_32b_x_32b(p1_array_index_58976, p1_array_index_58977);
  assign p2_smul_59364_comb = smul32b_32b_x_32b(p1_array_index_58978, p1_array_index_58979);
  assign p2_smul_59365_comb = smul32b_32b_x_32b(p1_array_index_58980, p1_array_index_58981);
  assign p2_smul_59366_comb = smul32b_32b_x_32b(p1_array_index_58982, p1_array_index_58983);
  assign p2_smul_59367_comb = smul32b_32b_x_32b(p1_array_index_58984, p1_array_index_58985);
  assign p2_smul_59368_comb = smul32b_32b_x_32b(p1_array_index_58986, p1_array_index_58987);
  assign p2_smul_59369_comb = smul32b_32b_x_32b(p1_array_index_58988, p1_array_index_58989);
  assign p2_add_60126_comb = p2_smul_59866_comb + p2_smul_59867_comb;
  assign p2_add_60127_comb = p2_smul_59868_comb + p2_smul_59869_comb;
  assign p2_add_60128_comb = p2_smul_59870_comb + p2_smul_59871_comb;
  assign p2_add_60129_comb = p2_smul_59872_comb + p2_smul_59873_comb;
  assign p2_add_60122_comb = p2_smul_59858_comb + p2_smul_59859_comb;
  assign p2_add_60123_comb = p2_smul_59860_comb + p2_smul_59861_comb;
  assign p2_add_60124_comb = p2_smul_59862_comb + p2_smul_59863_comb;
  assign p2_add_60125_comb = p2_smul_59864_comb + p2_smul_59865_comb;
  assign p2_add_60118_comb = p2_smul_59850_comb + p2_smul_59851_comb;
  assign p2_add_60119_comb = p2_smul_59852_comb + p2_smul_59853_comb;
  assign p2_add_60120_comb = p2_smul_59854_comb + p2_smul_59855_comb;
  assign p2_add_60121_comb = p2_smul_59856_comb + p2_smul_59857_comb;
  assign p2_add_60114_comb = p2_smul_59842_comb + p2_smul_59843_comb;
  assign p2_add_60115_comb = p2_smul_59844_comb + p2_smul_59845_comb;
  assign p2_add_60116_comb = p2_smul_59846_comb + p2_smul_59847_comb;
  assign p2_add_60117_comb = p2_smul_59848_comb + p2_smul_59849_comb;
  assign p2_add_60110_comb = p2_smul_59834_comb + p2_smul_59835_comb;
  assign p2_add_60111_comb = p2_smul_59836_comb + p2_smul_59837_comb;
  assign p2_add_60112_comb = p2_smul_59838_comb + p2_smul_59839_comb;
  assign p2_add_60113_comb = p2_smul_59840_comb + p2_smul_59841_comb;
  assign p2_add_60106_comb = p2_smul_59826_comb + p2_smul_59827_comb;
  assign p2_add_60107_comb = p2_smul_59828_comb + p2_smul_59829_comb;
  assign p2_add_60108_comb = p2_smul_59830_comb + p2_smul_59831_comb;
  assign p2_add_60109_comb = p2_smul_59832_comb + p2_smul_59833_comb;
  assign p2_add_60102_comb = p2_smul_59818_comb + p2_smul_59819_comb;
  assign p2_add_60103_comb = p2_smul_59820_comb + p2_smul_59821_comb;
  assign p2_add_60104_comb = p2_smul_59822_comb + p2_smul_59823_comb;
  assign p2_add_60105_comb = p2_smul_59824_comb + p2_smul_59825_comb;
  assign p2_add_60098_comb = p2_smul_59810_comb + p2_smul_59811_comb;
  assign p2_add_60099_comb = p2_smul_59812_comb + p2_smul_59813_comb;
  assign p2_add_60100_comb = p2_smul_59814_comb + p2_smul_59815_comb;
  assign p2_add_60101_comb = p2_smul_59816_comb + p2_smul_59817_comb;
  assign p2_add_60094_comb = p2_smul_59802_comb + p2_smul_59803_comb;
  assign p2_add_60095_comb = p2_smul_59804_comb + p2_smul_59805_comb;
  assign p2_add_60096_comb = p2_smul_59806_comb + p2_smul_59807_comb;
  assign p2_add_60097_comb = p2_smul_59808_comb + p2_smul_59809_comb;
  assign p2_add_60090_comb = p2_smul_59794_comb + p2_smul_59795_comb;
  assign p2_add_60091_comb = p2_smul_59796_comb + p2_smul_59797_comb;
  assign p2_add_60092_comb = p2_smul_59798_comb + p2_smul_59799_comb;
  assign p2_add_60093_comb = p2_smul_59800_comb + p2_smul_59801_comb;
  assign p2_add_60086_comb = p2_smul_59786_comb + p2_smul_59787_comb;
  assign p2_add_60087_comb = p2_smul_59788_comb + p2_smul_59789_comb;
  assign p2_add_60088_comb = p2_smul_59790_comb + p2_smul_59791_comb;
  assign p2_add_60089_comb = p2_smul_59792_comb + p2_smul_59793_comb;
  assign p2_add_60082_comb = p2_smul_59778_comb + p2_smul_59779_comb;
  assign p2_add_60083_comb = p2_smul_59780_comb + p2_smul_59781_comb;
  assign p2_add_60084_comb = p2_smul_59782_comb + p2_smul_59783_comb;
  assign p2_add_60085_comb = p2_smul_59784_comb + p2_smul_59785_comb;
  assign p2_add_60078_comb = p2_smul_59770_comb + p2_smul_59771_comb;
  assign p2_add_60079_comb = p2_smul_59772_comb + p2_smul_59773_comb;
  assign p2_add_60080_comb = p2_smul_59774_comb + p2_smul_59775_comb;
  assign p2_add_60081_comb = p2_smul_59776_comb + p2_smul_59777_comb;
  assign p2_add_60074_comb = p2_smul_59762_comb + p2_smul_59763_comb;
  assign p2_add_60075_comb = p2_smul_59764_comb + p2_smul_59765_comb;
  assign p2_add_60076_comb = p2_smul_59766_comb + p2_smul_59767_comb;
  assign p2_add_60077_comb = p2_smul_59768_comb + p2_smul_59769_comb;
  assign p2_add_60070_comb = p2_smul_59754_comb + p2_smul_59755_comb;
  assign p2_add_60071_comb = p2_smul_59756_comb + p2_smul_59757_comb;
  assign p2_add_60072_comb = p2_smul_59758_comb + p2_smul_59759_comb;
  assign p2_add_60073_comb = p2_smul_59760_comb + p2_smul_59761_comb;
  assign p2_add_60066_comb = p2_smul_59746_comb + p2_smul_59747_comb;
  assign p2_add_60067_comb = p2_smul_59748_comb + p2_smul_59749_comb;
  assign p2_add_60068_comb = p2_smul_59750_comb + p2_smul_59751_comb;
  assign p2_add_60069_comb = p2_smul_59752_comb + p2_smul_59753_comb;
  assign p2_add_60062_comb = p2_smul_59738_comb + p2_smul_59739_comb;
  assign p2_add_60063_comb = p2_smul_59740_comb + p2_smul_59741_comb;
  assign p2_add_60064_comb = p2_smul_59742_comb + p2_smul_59743_comb;
  assign p2_add_60065_comb = p2_smul_59744_comb + p2_smul_59745_comb;
  assign p2_add_60058_comb = p2_smul_59730_comb + p2_smul_59731_comb;
  assign p2_add_60059_comb = p2_smul_59732_comb + p2_smul_59733_comb;
  assign p2_add_60060_comb = p2_smul_59734_comb + p2_smul_59735_comb;
  assign p2_add_60061_comb = p2_smul_59736_comb + p2_smul_59737_comb;
  assign p2_add_60054_comb = p2_smul_59722_comb + p2_smul_59723_comb;
  assign p2_add_60055_comb = p2_smul_59724_comb + p2_smul_59725_comb;
  assign p2_add_60056_comb = p2_smul_59726_comb + p2_smul_59727_comb;
  assign p2_add_60057_comb = p2_smul_59728_comb + p2_smul_59729_comb;
  assign p2_add_60050_comb = p2_smul_59714_comb + p2_smul_59715_comb;
  assign p2_add_60051_comb = p2_smul_59716_comb + p2_smul_59717_comb;
  assign p2_add_60052_comb = p2_smul_59718_comb + p2_smul_59719_comb;
  assign p2_add_60053_comb = p2_smul_59720_comb + p2_smul_59721_comb;
  assign p2_add_60046_comb = p2_smul_59706_comb + p2_smul_59707_comb;
  assign p2_add_60047_comb = p2_smul_59708_comb + p2_smul_59709_comb;
  assign p2_add_60048_comb = p2_smul_59710_comb + p2_smul_59711_comb;
  assign p2_add_60049_comb = p2_smul_59712_comb + p2_smul_59713_comb;
  assign p2_add_60042_comb = p2_smul_59698_comb + p2_smul_59699_comb;
  assign p2_add_60043_comb = p2_smul_59700_comb + p2_smul_59701_comb;
  assign p2_add_60044_comb = p2_smul_59702_comb + p2_smul_59703_comb;
  assign p2_add_60045_comb = p2_smul_59704_comb + p2_smul_59705_comb;
  assign p2_add_60038_comb = p2_smul_59690_comb + p2_smul_59691_comb;
  assign p2_add_60039_comb = p2_smul_59692_comb + p2_smul_59693_comb;
  assign p2_add_60040_comb = p2_smul_59694_comb + p2_smul_59695_comb;
  assign p2_add_60041_comb = p2_smul_59696_comb + p2_smul_59697_comb;
  assign p2_add_60034_comb = p2_smul_59682_comb + p2_smul_59683_comb;
  assign p2_add_60035_comb = p2_smul_59684_comb + p2_smul_59685_comb;
  assign p2_add_60036_comb = p2_smul_59686_comb + p2_smul_59687_comb;
  assign p2_add_60037_comb = p2_smul_59688_comb + p2_smul_59689_comb;
  assign p2_add_60030_comb = p2_smul_59674_comb + p2_smul_59675_comb;
  assign p2_add_60031_comb = p2_smul_59676_comb + p2_smul_59677_comb;
  assign p2_add_60032_comb = p2_smul_59678_comb + p2_smul_59679_comb;
  assign p2_add_60033_comb = p2_smul_59680_comb + p2_smul_59681_comb;
  assign p2_add_60026_comb = p2_smul_59666_comb + p2_smul_59667_comb;
  assign p2_add_60027_comb = p2_smul_59668_comb + p2_smul_59669_comb;
  assign p2_add_60028_comb = p2_smul_59670_comb + p2_smul_59671_comb;
  assign p2_add_60029_comb = p2_smul_59672_comb + p2_smul_59673_comb;
  assign p2_add_60022_comb = p2_smul_59658_comb + p2_smul_59659_comb;
  assign p2_add_60023_comb = p2_smul_59660_comb + p2_smul_59661_comb;
  assign p2_add_60024_comb = p2_smul_59662_comb + p2_smul_59663_comb;
  assign p2_add_60025_comb = p2_smul_59664_comb + p2_smul_59665_comb;
  assign p2_add_60018_comb = p2_smul_59650_comb + p2_smul_59651_comb;
  assign p2_add_60019_comb = p2_smul_59652_comb + p2_smul_59653_comb;
  assign p2_add_60020_comb = p2_smul_59654_comb + p2_smul_59655_comb;
  assign p2_add_60021_comb = p2_smul_59656_comb + p2_smul_59657_comb;
  assign p2_add_60014_comb = p2_smul_59642_comb + p2_smul_59643_comb;
  assign p2_add_60015_comb = p2_smul_59644_comb + p2_smul_59645_comb;
  assign p2_add_60016_comb = p2_smul_59646_comb + p2_smul_59647_comb;
  assign p2_add_60017_comb = p2_smul_59648_comb + p2_smul_59649_comb;
  assign p2_add_60010_comb = p2_smul_59634_comb + p2_smul_59635_comb;
  assign p2_add_60011_comb = p2_smul_59636_comb + p2_smul_59637_comb;
  assign p2_add_60012_comb = p2_smul_59638_comb + p2_smul_59639_comb;
  assign p2_add_60013_comb = p2_smul_59640_comb + p2_smul_59641_comb;
  assign p2_add_60006_comb = p2_smul_59626_comb + p2_smul_59627_comb;
  assign p2_add_60007_comb = p2_smul_59628_comb + p2_smul_59629_comb;
  assign p2_add_60008_comb = p2_smul_59630_comb + p2_smul_59631_comb;
  assign p2_add_60009_comb = p2_smul_59632_comb + p2_smul_59633_comb;
  assign p2_add_60002_comb = p2_smul_59618_comb + p2_smul_59619_comb;
  assign p2_add_60003_comb = p2_smul_59620_comb + p2_smul_59621_comb;
  assign p2_add_60004_comb = p2_smul_59622_comb + p2_smul_59623_comb;
  assign p2_add_60005_comb = p2_smul_59624_comb + p2_smul_59625_comb;
  assign p2_add_59998_comb = p2_smul_59610_comb + p2_smul_59611_comb;
  assign p2_add_59999_comb = p2_smul_59612_comb + p2_smul_59613_comb;
  assign p2_add_60000_comb = p2_smul_59614_comb + p2_smul_59615_comb;
  assign p2_add_60001_comb = p2_smul_59616_comb + p2_smul_59617_comb;
  assign p2_add_59994_comb = p2_smul_59602_comb + p2_smul_59603_comb;
  assign p2_add_59995_comb = p2_smul_59604_comb + p2_smul_59605_comb;
  assign p2_add_59996_comb = p2_smul_59606_comb + p2_smul_59607_comb;
  assign p2_add_59997_comb = p2_smul_59608_comb + p2_smul_59609_comb;
  assign p2_add_59990_comb = p2_smul_59594_comb + p2_smul_59595_comb;
  assign p2_add_59991_comb = p2_smul_59596_comb + p2_smul_59597_comb;
  assign p2_add_59992_comb = p2_smul_59598_comb + p2_smul_59599_comb;
  assign p2_add_59993_comb = p2_smul_59600_comb + p2_smul_59601_comb;
  assign p2_add_59986_comb = p2_smul_59586_comb + p2_smul_59587_comb;
  assign p2_add_59987_comb = p2_smul_59588_comb + p2_smul_59589_comb;
  assign p2_add_59988_comb = p2_smul_59590_comb + p2_smul_59591_comb;
  assign p2_add_59989_comb = p2_smul_59592_comb + p2_smul_59593_comb;
  assign p2_add_59982_comb = p2_smul_59578_comb + p2_smul_59579_comb;
  assign p2_add_59983_comb = p2_smul_59580_comb + p2_smul_59581_comb;
  assign p2_add_59984_comb = p2_smul_59582_comb + p2_smul_59583_comb;
  assign p2_add_59985_comb = p2_smul_59584_comb + p2_smul_59585_comb;
  assign p2_add_59978_comb = p2_smul_59570_comb + p2_smul_59571_comb;
  assign p2_add_59979_comb = p2_smul_59572_comb + p2_smul_59573_comb;
  assign p2_add_59980_comb = p2_smul_59574_comb + p2_smul_59575_comb;
  assign p2_add_59981_comb = p2_smul_59576_comb + p2_smul_59577_comb;
  assign p2_add_59974_comb = p2_smul_59562_comb + p2_smul_59563_comb;
  assign p2_add_59975_comb = p2_smul_59564_comb + p2_smul_59565_comb;
  assign p2_add_59976_comb = p2_smul_59566_comb + p2_smul_59567_comb;
  assign p2_add_59977_comb = p2_smul_59568_comb + p2_smul_59569_comb;
  assign p2_add_59970_comb = p2_smul_59554_comb + p2_smul_59555_comb;
  assign p2_add_59971_comb = p2_smul_59556_comb + p2_smul_59557_comb;
  assign p2_add_59972_comb = p2_smul_59558_comb + p2_smul_59559_comb;
  assign p2_add_59973_comb = p2_smul_59560_comb + p2_smul_59561_comb;
  assign p2_add_59966_comb = p2_smul_59546_comb + p2_smul_59547_comb;
  assign p2_add_59967_comb = p2_smul_59548_comb + p2_smul_59549_comb;
  assign p2_add_59968_comb = p2_smul_59550_comb + p2_smul_59551_comb;
  assign p2_add_59969_comb = p2_smul_59552_comb + p2_smul_59553_comb;
  assign p2_add_59962_comb = p2_smul_59538_comb + p2_smul_59539_comb;
  assign p2_add_59963_comb = p2_smul_59540_comb + p2_smul_59541_comb;
  assign p2_add_59964_comb = p2_smul_59542_comb + p2_smul_59543_comb;
  assign p2_add_59965_comb = p2_smul_59544_comb + p2_smul_59545_comb;
  assign p2_add_59958_comb = p2_smul_59530_comb + p2_smul_59531_comb;
  assign p2_add_59959_comb = p2_smul_59532_comb + p2_smul_59533_comb;
  assign p2_add_59960_comb = p2_smul_59534_comb + p2_smul_59535_comb;
  assign p2_add_59961_comb = p2_smul_59536_comb + p2_smul_59537_comb;
  assign p2_add_59954_comb = p2_smul_59522_comb + p2_smul_59523_comb;
  assign p2_add_59955_comb = p2_smul_59524_comb + p2_smul_59525_comb;
  assign p2_add_59956_comb = p2_smul_59526_comb + p2_smul_59527_comb;
  assign p2_add_59957_comb = p2_smul_59528_comb + p2_smul_59529_comb;
  assign p2_add_59950_comb = p2_smul_59514_comb + p2_smul_59515_comb;
  assign p2_add_59951_comb = p2_smul_59516_comb + p2_smul_59517_comb;
  assign p2_add_59952_comb = p2_smul_59518_comb + p2_smul_59519_comb;
  assign p2_add_59953_comb = p2_smul_59520_comb + p2_smul_59521_comb;
  assign p2_add_59946_comb = p2_smul_59506_comb + p2_smul_59507_comb;
  assign p2_add_59947_comb = p2_smul_59508_comb + p2_smul_59509_comb;
  assign p2_add_59948_comb = p2_smul_59510_comb + p2_smul_59511_comb;
  assign p2_add_59949_comb = p2_smul_59512_comb + p2_smul_59513_comb;
  assign p2_add_59942_comb = p2_smul_59498_comb + p2_smul_59499_comb;
  assign p2_add_59943_comb = p2_smul_59500_comb + p2_smul_59501_comb;
  assign p2_add_59944_comb = p2_smul_59502_comb + p2_smul_59503_comb;
  assign p2_add_59945_comb = p2_smul_59504_comb + p2_smul_59505_comb;
  assign p2_add_59938_comb = p2_smul_59490_comb + p2_smul_59491_comb;
  assign p2_add_59939_comb = p2_smul_59492_comb + p2_smul_59493_comb;
  assign p2_add_59940_comb = p2_smul_59494_comb + p2_smul_59495_comb;
  assign p2_add_59941_comb = p2_smul_59496_comb + p2_smul_59497_comb;
  assign p2_add_59934_comb = p2_smul_59482_comb + p2_smul_59483_comb;
  assign p2_add_59935_comb = p2_smul_59484_comb + p2_smul_59485_comb;
  assign p2_add_59936_comb = p2_smul_59486_comb + p2_smul_59487_comb;
  assign p2_add_59937_comb = p2_smul_59488_comb + p2_smul_59489_comb;
  assign p2_add_59930_comb = p2_smul_59474_comb + p2_smul_59475_comb;
  assign p2_add_59931_comb = p2_smul_59476_comb + p2_smul_59477_comb;
  assign p2_add_59932_comb = p2_smul_59478_comb + p2_smul_59479_comb;
  assign p2_add_59933_comb = p2_smul_59480_comb + p2_smul_59481_comb;
  assign p2_add_59926_comb = p2_smul_59466_comb + p2_smul_59467_comb;
  assign p2_add_59927_comb = p2_smul_59468_comb + p2_smul_59469_comb;
  assign p2_add_59928_comb = p2_smul_59470_comb + p2_smul_59471_comb;
  assign p2_add_59929_comb = p2_smul_59472_comb + p2_smul_59473_comb;
  assign p2_add_59922_comb = p2_smul_59458_comb + p2_smul_59459_comb;
  assign p2_add_59923_comb = p2_smul_59460_comb + p2_smul_59461_comb;
  assign p2_add_59924_comb = p2_smul_59462_comb + p2_smul_59463_comb;
  assign p2_add_59925_comb = p2_smul_59464_comb + p2_smul_59465_comb;
  assign p2_add_59918_comb = p2_smul_59450_comb + p2_smul_59451_comb;
  assign p2_add_59919_comb = p2_smul_59452_comb + p2_smul_59453_comb;
  assign p2_add_59920_comb = p2_smul_59454_comb + p2_smul_59455_comb;
  assign p2_add_59921_comb = p2_smul_59456_comb + p2_smul_59457_comb;
  assign p2_add_59914_comb = p2_smul_59442_comb + p2_smul_59443_comb;
  assign p2_add_59915_comb = p2_smul_59444_comb + p2_smul_59445_comb;
  assign p2_add_59916_comb = p2_smul_59446_comb + p2_smul_59447_comb;
  assign p2_add_59917_comb = p2_smul_59448_comb + p2_smul_59449_comb;
  assign p2_add_59910_comb = p2_smul_59434_comb + p2_smul_59435_comb;
  assign p2_add_59911_comb = p2_smul_59436_comb + p2_smul_59437_comb;
  assign p2_add_59912_comb = p2_smul_59438_comb + p2_smul_59439_comb;
  assign p2_add_59913_comb = p2_smul_59440_comb + p2_smul_59441_comb;
  assign p2_add_59906_comb = p2_smul_59426_comb + p2_smul_59427_comb;
  assign p2_add_59907_comb = p2_smul_59428_comb + p2_smul_59429_comb;
  assign p2_add_59908_comb = p2_smul_59430_comb + p2_smul_59431_comb;
  assign p2_add_59909_comb = p2_smul_59432_comb + p2_smul_59433_comb;
  assign p2_add_59902_comb = p2_smul_59418_comb + p2_smul_59419_comb;
  assign p2_add_59903_comb = p2_smul_59420_comb + p2_smul_59421_comb;
  assign p2_add_59904_comb = p2_smul_59422_comb + p2_smul_59423_comb;
  assign p2_add_59905_comb = p2_smul_59424_comb + p2_smul_59425_comb;
  assign p2_add_59898_comb = p2_smul_59410_comb + p2_smul_59411_comb;
  assign p2_add_59899_comb = p2_smul_59412_comb + p2_smul_59413_comb;
  assign p2_add_59900_comb = p2_smul_59414_comb + p2_smul_59415_comb;
  assign p2_add_59901_comb = p2_smul_59416_comb + p2_smul_59417_comb;
  assign p2_add_59894_comb = p2_smul_59402_comb + p2_smul_59403_comb;
  assign p2_add_59895_comb = p2_smul_59404_comb + p2_smul_59405_comb;
  assign p2_add_59896_comb = p2_smul_59406_comb + p2_smul_59407_comb;
  assign p2_add_59897_comb = p2_smul_59408_comb + p2_smul_59409_comb;
  assign p2_add_59890_comb = p2_smul_59394_comb + p2_smul_59395_comb;
  assign p2_add_59891_comb = p2_smul_59396_comb + p2_smul_59397_comb;
  assign p2_add_59892_comb = p2_smul_59398_comb + p2_smul_59399_comb;
  assign p2_add_59893_comb = p2_smul_59400_comb + p2_smul_59401_comb;
  assign p2_add_59886_comb = p2_smul_59386_comb + p2_smul_59387_comb;
  assign p2_add_59887_comb = p2_smul_59388_comb + p2_smul_59389_comb;
  assign p2_add_59888_comb = p2_smul_59390_comb + p2_smul_59391_comb;
  assign p2_add_59889_comb = p2_smul_59392_comb + p2_smul_59393_comb;
  assign p2_add_59882_comb = p2_smul_59378_comb + p2_smul_59379_comb;
  assign p2_add_59883_comb = p2_smul_59380_comb + p2_smul_59381_comb;
  assign p2_add_59884_comb = p2_smul_59382_comb + p2_smul_59383_comb;
  assign p2_add_59885_comb = p2_smul_59384_comb + p2_smul_59385_comb;
  assign p2_add_59878_comb = p2_smul_59370_comb + p2_smul_59371_comb;
  assign p2_add_59879_comb = p2_smul_59372_comb + p2_smul_59373_comb;
  assign p2_add_59880_comb = p2_smul_59374_comb + p2_smul_59375_comb;
  assign p2_add_59881_comb = p2_smul_59376_comb + p2_smul_59377_comb;
  assign p2_add_59874_comb = p2_smul_59362_comb + p2_smul_59363_comb;
  assign p2_add_59875_comb = p2_smul_59364_comb + p2_smul_59365_comb;
  assign p2_add_59876_comb = p2_smul_59366_comb + p2_smul_59367_comb;
  assign p2_add_59877_comb = p2_smul_59368_comb + p2_smul_59369_comb;

  // Registers for pipe stage 2:
  reg [31:0] p2_a[8][8];
  reg [31:0] p2_b[8][8];
  reg [31:0] p2_add_60126;
  reg [31:0] p2_add_60127;
  reg [31:0] p2_add_60128;
  reg [31:0] p2_add_60129;
  reg [31:0] p2_add_60122;
  reg [31:0] p2_add_60123;
  reg [31:0] p2_add_60124;
  reg [31:0] p2_add_60125;
  reg [31:0] p2_add_60118;
  reg [31:0] p2_add_60119;
  reg [31:0] p2_add_60120;
  reg [31:0] p2_add_60121;
  reg [31:0] p2_add_60114;
  reg [31:0] p2_add_60115;
  reg [31:0] p2_add_60116;
  reg [31:0] p2_add_60117;
  reg [31:0] p2_add_60110;
  reg [31:0] p2_add_60111;
  reg [31:0] p2_add_60112;
  reg [31:0] p2_add_60113;
  reg [31:0] p2_add_60106;
  reg [31:0] p2_add_60107;
  reg [31:0] p2_add_60108;
  reg [31:0] p2_add_60109;
  reg [31:0] p2_add_60102;
  reg [31:0] p2_add_60103;
  reg [31:0] p2_add_60104;
  reg [31:0] p2_add_60105;
  reg [31:0] p2_add_60098;
  reg [31:0] p2_add_60099;
  reg [31:0] p2_add_60100;
  reg [31:0] p2_add_60101;
  reg [31:0] p2_add_60094;
  reg [31:0] p2_add_60095;
  reg [31:0] p2_add_60096;
  reg [31:0] p2_add_60097;
  reg [31:0] p2_add_60090;
  reg [31:0] p2_add_60091;
  reg [31:0] p2_add_60092;
  reg [31:0] p2_add_60093;
  reg [31:0] p2_add_60086;
  reg [31:0] p2_add_60087;
  reg [31:0] p2_add_60088;
  reg [31:0] p2_add_60089;
  reg [31:0] p2_add_60082;
  reg [31:0] p2_add_60083;
  reg [31:0] p2_add_60084;
  reg [31:0] p2_add_60085;
  reg [31:0] p2_add_60078;
  reg [31:0] p2_add_60079;
  reg [31:0] p2_add_60080;
  reg [31:0] p2_add_60081;
  reg [31:0] p2_add_60074;
  reg [31:0] p2_add_60075;
  reg [31:0] p2_add_60076;
  reg [31:0] p2_add_60077;
  reg [31:0] p2_add_60070;
  reg [31:0] p2_add_60071;
  reg [31:0] p2_add_60072;
  reg [31:0] p2_add_60073;
  reg [31:0] p2_add_60066;
  reg [31:0] p2_add_60067;
  reg [31:0] p2_add_60068;
  reg [31:0] p2_add_60069;
  reg [31:0] p2_add_60062;
  reg [31:0] p2_add_60063;
  reg [31:0] p2_add_60064;
  reg [31:0] p2_add_60065;
  reg [31:0] p2_add_60058;
  reg [31:0] p2_add_60059;
  reg [31:0] p2_add_60060;
  reg [31:0] p2_add_60061;
  reg [31:0] p2_add_60054;
  reg [31:0] p2_add_60055;
  reg [31:0] p2_add_60056;
  reg [31:0] p2_add_60057;
  reg [31:0] p2_add_60050;
  reg [31:0] p2_add_60051;
  reg [31:0] p2_add_60052;
  reg [31:0] p2_add_60053;
  reg [31:0] p2_add_60046;
  reg [31:0] p2_add_60047;
  reg [31:0] p2_add_60048;
  reg [31:0] p2_add_60049;
  reg [31:0] p2_add_60042;
  reg [31:0] p2_add_60043;
  reg [31:0] p2_add_60044;
  reg [31:0] p2_add_60045;
  reg [31:0] p2_add_60038;
  reg [31:0] p2_add_60039;
  reg [31:0] p2_add_60040;
  reg [31:0] p2_add_60041;
  reg [31:0] p2_add_60034;
  reg [31:0] p2_add_60035;
  reg [31:0] p2_add_60036;
  reg [31:0] p2_add_60037;
  reg [31:0] p2_add_60030;
  reg [31:0] p2_add_60031;
  reg [31:0] p2_add_60032;
  reg [31:0] p2_add_60033;
  reg [31:0] p2_add_60026;
  reg [31:0] p2_add_60027;
  reg [31:0] p2_add_60028;
  reg [31:0] p2_add_60029;
  reg [31:0] p2_add_60022;
  reg [31:0] p2_add_60023;
  reg [31:0] p2_add_60024;
  reg [31:0] p2_add_60025;
  reg [31:0] p2_add_60018;
  reg [31:0] p2_add_60019;
  reg [31:0] p2_add_60020;
  reg [31:0] p2_add_60021;
  reg [31:0] p2_add_60014;
  reg [31:0] p2_add_60015;
  reg [31:0] p2_add_60016;
  reg [31:0] p2_add_60017;
  reg [31:0] p2_add_60010;
  reg [31:0] p2_add_60011;
  reg [31:0] p2_add_60012;
  reg [31:0] p2_add_60013;
  reg [31:0] p2_add_60006;
  reg [31:0] p2_add_60007;
  reg [31:0] p2_add_60008;
  reg [31:0] p2_add_60009;
  reg [31:0] p2_add_60002;
  reg [31:0] p2_add_60003;
  reg [31:0] p2_add_60004;
  reg [31:0] p2_add_60005;
  reg [31:0] p2_add_59998;
  reg [31:0] p2_add_59999;
  reg [31:0] p2_add_60000;
  reg [31:0] p2_add_60001;
  reg [31:0] p2_add_59994;
  reg [31:0] p2_add_59995;
  reg [31:0] p2_add_59996;
  reg [31:0] p2_add_59997;
  reg [31:0] p2_add_59990;
  reg [31:0] p2_add_59991;
  reg [31:0] p2_add_59992;
  reg [31:0] p2_add_59993;
  reg [31:0] p2_add_59986;
  reg [31:0] p2_add_59987;
  reg [31:0] p2_add_59988;
  reg [31:0] p2_add_59989;
  reg [31:0] p2_add_59982;
  reg [31:0] p2_add_59983;
  reg [31:0] p2_add_59984;
  reg [31:0] p2_add_59985;
  reg [31:0] p2_add_59978;
  reg [31:0] p2_add_59979;
  reg [31:0] p2_add_59980;
  reg [31:0] p2_add_59981;
  reg [31:0] p2_add_59974;
  reg [31:0] p2_add_59975;
  reg [31:0] p2_add_59976;
  reg [31:0] p2_add_59977;
  reg [31:0] p2_add_59970;
  reg [31:0] p2_add_59971;
  reg [31:0] p2_add_59972;
  reg [31:0] p2_add_59973;
  reg [31:0] p2_add_59966;
  reg [31:0] p2_add_59967;
  reg [31:0] p2_add_59968;
  reg [31:0] p2_add_59969;
  reg [31:0] p2_add_59962;
  reg [31:0] p2_add_59963;
  reg [31:0] p2_add_59964;
  reg [31:0] p2_add_59965;
  reg [31:0] p2_add_59958;
  reg [31:0] p2_add_59959;
  reg [31:0] p2_add_59960;
  reg [31:0] p2_add_59961;
  reg [31:0] p2_add_59954;
  reg [31:0] p2_add_59955;
  reg [31:0] p2_add_59956;
  reg [31:0] p2_add_59957;
  reg [31:0] p2_add_59950;
  reg [31:0] p2_add_59951;
  reg [31:0] p2_add_59952;
  reg [31:0] p2_add_59953;
  reg [31:0] p2_add_59946;
  reg [31:0] p2_add_59947;
  reg [31:0] p2_add_59948;
  reg [31:0] p2_add_59949;
  reg [31:0] p2_add_59942;
  reg [31:0] p2_add_59943;
  reg [31:0] p2_add_59944;
  reg [31:0] p2_add_59945;
  reg [31:0] p2_add_59938;
  reg [31:0] p2_add_59939;
  reg [31:0] p2_add_59940;
  reg [31:0] p2_add_59941;
  reg [31:0] p2_add_59934;
  reg [31:0] p2_add_59935;
  reg [31:0] p2_add_59936;
  reg [31:0] p2_add_59937;
  reg [31:0] p2_add_59930;
  reg [31:0] p2_add_59931;
  reg [31:0] p2_add_59932;
  reg [31:0] p2_add_59933;
  reg [31:0] p2_add_59926;
  reg [31:0] p2_add_59927;
  reg [31:0] p2_add_59928;
  reg [31:0] p2_add_59929;
  reg [31:0] p2_add_59922;
  reg [31:0] p2_add_59923;
  reg [31:0] p2_add_59924;
  reg [31:0] p2_add_59925;
  reg [31:0] p2_add_59918;
  reg [31:0] p2_add_59919;
  reg [31:0] p2_add_59920;
  reg [31:0] p2_add_59921;
  reg [31:0] p2_add_59914;
  reg [31:0] p2_add_59915;
  reg [31:0] p2_add_59916;
  reg [31:0] p2_add_59917;
  reg [31:0] p2_add_59910;
  reg [31:0] p2_add_59911;
  reg [31:0] p2_add_59912;
  reg [31:0] p2_add_59913;
  reg [31:0] p2_add_59906;
  reg [31:0] p2_add_59907;
  reg [31:0] p2_add_59908;
  reg [31:0] p2_add_59909;
  reg [31:0] p2_add_59902;
  reg [31:0] p2_add_59903;
  reg [31:0] p2_add_59904;
  reg [31:0] p2_add_59905;
  reg [31:0] p2_add_59898;
  reg [31:0] p2_add_59899;
  reg [31:0] p2_add_59900;
  reg [31:0] p2_add_59901;
  reg [31:0] p2_add_59894;
  reg [31:0] p2_add_59895;
  reg [31:0] p2_add_59896;
  reg [31:0] p2_add_59897;
  reg [31:0] p2_add_59890;
  reg [31:0] p2_add_59891;
  reg [31:0] p2_add_59892;
  reg [31:0] p2_add_59893;
  reg [31:0] p2_add_59886;
  reg [31:0] p2_add_59887;
  reg [31:0] p2_add_59888;
  reg [31:0] p2_add_59889;
  reg [31:0] p2_add_59882;
  reg [31:0] p2_add_59883;
  reg [31:0] p2_add_59884;
  reg [31:0] p2_add_59885;
  reg [31:0] p2_add_59878;
  reg [31:0] p2_add_59879;
  reg [31:0] p2_add_59880;
  reg [31:0] p2_add_59881;
  reg [31:0] p2_add_59874;
  reg [31:0] p2_add_59875;
  reg [31:0] p2_add_59876;
  reg [31:0] p2_add_59877;
  always_ff @ (posedge clk) begin
    p2_a <= p1_a;
    p2_b <= p1_b;
    p2_add_60126 <= p2_add_60126_comb;
    p2_add_60127 <= p2_add_60127_comb;
    p2_add_60128 <= p2_add_60128_comb;
    p2_add_60129 <= p2_add_60129_comb;
    p2_add_60122 <= p2_add_60122_comb;
    p2_add_60123 <= p2_add_60123_comb;
    p2_add_60124 <= p2_add_60124_comb;
    p2_add_60125 <= p2_add_60125_comb;
    p2_add_60118 <= p2_add_60118_comb;
    p2_add_60119 <= p2_add_60119_comb;
    p2_add_60120 <= p2_add_60120_comb;
    p2_add_60121 <= p2_add_60121_comb;
    p2_add_60114 <= p2_add_60114_comb;
    p2_add_60115 <= p2_add_60115_comb;
    p2_add_60116 <= p2_add_60116_comb;
    p2_add_60117 <= p2_add_60117_comb;
    p2_add_60110 <= p2_add_60110_comb;
    p2_add_60111 <= p2_add_60111_comb;
    p2_add_60112 <= p2_add_60112_comb;
    p2_add_60113 <= p2_add_60113_comb;
    p2_add_60106 <= p2_add_60106_comb;
    p2_add_60107 <= p2_add_60107_comb;
    p2_add_60108 <= p2_add_60108_comb;
    p2_add_60109 <= p2_add_60109_comb;
    p2_add_60102 <= p2_add_60102_comb;
    p2_add_60103 <= p2_add_60103_comb;
    p2_add_60104 <= p2_add_60104_comb;
    p2_add_60105 <= p2_add_60105_comb;
    p2_add_60098 <= p2_add_60098_comb;
    p2_add_60099 <= p2_add_60099_comb;
    p2_add_60100 <= p2_add_60100_comb;
    p2_add_60101 <= p2_add_60101_comb;
    p2_add_60094 <= p2_add_60094_comb;
    p2_add_60095 <= p2_add_60095_comb;
    p2_add_60096 <= p2_add_60096_comb;
    p2_add_60097 <= p2_add_60097_comb;
    p2_add_60090 <= p2_add_60090_comb;
    p2_add_60091 <= p2_add_60091_comb;
    p2_add_60092 <= p2_add_60092_comb;
    p2_add_60093 <= p2_add_60093_comb;
    p2_add_60086 <= p2_add_60086_comb;
    p2_add_60087 <= p2_add_60087_comb;
    p2_add_60088 <= p2_add_60088_comb;
    p2_add_60089 <= p2_add_60089_comb;
    p2_add_60082 <= p2_add_60082_comb;
    p2_add_60083 <= p2_add_60083_comb;
    p2_add_60084 <= p2_add_60084_comb;
    p2_add_60085 <= p2_add_60085_comb;
    p2_add_60078 <= p2_add_60078_comb;
    p2_add_60079 <= p2_add_60079_comb;
    p2_add_60080 <= p2_add_60080_comb;
    p2_add_60081 <= p2_add_60081_comb;
    p2_add_60074 <= p2_add_60074_comb;
    p2_add_60075 <= p2_add_60075_comb;
    p2_add_60076 <= p2_add_60076_comb;
    p2_add_60077 <= p2_add_60077_comb;
    p2_add_60070 <= p2_add_60070_comb;
    p2_add_60071 <= p2_add_60071_comb;
    p2_add_60072 <= p2_add_60072_comb;
    p2_add_60073 <= p2_add_60073_comb;
    p2_add_60066 <= p2_add_60066_comb;
    p2_add_60067 <= p2_add_60067_comb;
    p2_add_60068 <= p2_add_60068_comb;
    p2_add_60069 <= p2_add_60069_comb;
    p2_add_60062 <= p2_add_60062_comb;
    p2_add_60063 <= p2_add_60063_comb;
    p2_add_60064 <= p2_add_60064_comb;
    p2_add_60065 <= p2_add_60065_comb;
    p2_add_60058 <= p2_add_60058_comb;
    p2_add_60059 <= p2_add_60059_comb;
    p2_add_60060 <= p2_add_60060_comb;
    p2_add_60061 <= p2_add_60061_comb;
    p2_add_60054 <= p2_add_60054_comb;
    p2_add_60055 <= p2_add_60055_comb;
    p2_add_60056 <= p2_add_60056_comb;
    p2_add_60057 <= p2_add_60057_comb;
    p2_add_60050 <= p2_add_60050_comb;
    p2_add_60051 <= p2_add_60051_comb;
    p2_add_60052 <= p2_add_60052_comb;
    p2_add_60053 <= p2_add_60053_comb;
    p2_add_60046 <= p2_add_60046_comb;
    p2_add_60047 <= p2_add_60047_comb;
    p2_add_60048 <= p2_add_60048_comb;
    p2_add_60049 <= p2_add_60049_comb;
    p2_add_60042 <= p2_add_60042_comb;
    p2_add_60043 <= p2_add_60043_comb;
    p2_add_60044 <= p2_add_60044_comb;
    p2_add_60045 <= p2_add_60045_comb;
    p2_add_60038 <= p2_add_60038_comb;
    p2_add_60039 <= p2_add_60039_comb;
    p2_add_60040 <= p2_add_60040_comb;
    p2_add_60041 <= p2_add_60041_comb;
    p2_add_60034 <= p2_add_60034_comb;
    p2_add_60035 <= p2_add_60035_comb;
    p2_add_60036 <= p2_add_60036_comb;
    p2_add_60037 <= p2_add_60037_comb;
    p2_add_60030 <= p2_add_60030_comb;
    p2_add_60031 <= p2_add_60031_comb;
    p2_add_60032 <= p2_add_60032_comb;
    p2_add_60033 <= p2_add_60033_comb;
    p2_add_60026 <= p2_add_60026_comb;
    p2_add_60027 <= p2_add_60027_comb;
    p2_add_60028 <= p2_add_60028_comb;
    p2_add_60029 <= p2_add_60029_comb;
    p2_add_60022 <= p2_add_60022_comb;
    p2_add_60023 <= p2_add_60023_comb;
    p2_add_60024 <= p2_add_60024_comb;
    p2_add_60025 <= p2_add_60025_comb;
    p2_add_60018 <= p2_add_60018_comb;
    p2_add_60019 <= p2_add_60019_comb;
    p2_add_60020 <= p2_add_60020_comb;
    p2_add_60021 <= p2_add_60021_comb;
    p2_add_60014 <= p2_add_60014_comb;
    p2_add_60015 <= p2_add_60015_comb;
    p2_add_60016 <= p2_add_60016_comb;
    p2_add_60017 <= p2_add_60017_comb;
    p2_add_60010 <= p2_add_60010_comb;
    p2_add_60011 <= p2_add_60011_comb;
    p2_add_60012 <= p2_add_60012_comb;
    p2_add_60013 <= p2_add_60013_comb;
    p2_add_60006 <= p2_add_60006_comb;
    p2_add_60007 <= p2_add_60007_comb;
    p2_add_60008 <= p2_add_60008_comb;
    p2_add_60009 <= p2_add_60009_comb;
    p2_add_60002 <= p2_add_60002_comb;
    p2_add_60003 <= p2_add_60003_comb;
    p2_add_60004 <= p2_add_60004_comb;
    p2_add_60005 <= p2_add_60005_comb;
    p2_add_59998 <= p2_add_59998_comb;
    p2_add_59999 <= p2_add_59999_comb;
    p2_add_60000 <= p2_add_60000_comb;
    p2_add_60001 <= p2_add_60001_comb;
    p2_add_59994 <= p2_add_59994_comb;
    p2_add_59995 <= p2_add_59995_comb;
    p2_add_59996 <= p2_add_59996_comb;
    p2_add_59997 <= p2_add_59997_comb;
    p2_add_59990 <= p2_add_59990_comb;
    p2_add_59991 <= p2_add_59991_comb;
    p2_add_59992 <= p2_add_59992_comb;
    p2_add_59993 <= p2_add_59993_comb;
    p2_add_59986 <= p2_add_59986_comb;
    p2_add_59987 <= p2_add_59987_comb;
    p2_add_59988 <= p2_add_59988_comb;
    p2_add_59989 <= p2_add_59989_comb;
    p2_add_59982 <= p2_add_59982_comb;
    p2_add_59983 <= p2_add_59983_comb;
    p2_add_59984 <= p2_add_59984_comb;
    p2_add_59985 <= p2_add_59985_comb;
    p2_add_59978 <= p2_add_59978_comb;
    p2_add_59979 <= p2_add_59979_comb;
    p2_add_59980 <= p2_add_59980_comb;
    p2_add_59981 <= p2_add_59981_comb;
    p2_add_59974 <= p2_add_59974_comb;
    p2_add_59975 <= p2_add_59975_comb;
    p2_add_59976 <= p2_add_59976_comb;
    p2_add_59977 <= p2_add_59977_comb;
    p2_add_59970 <= p2_add_59970_comb;
    p2_add_59971 <= p2_add_59971_comb;
    p2_add_59972 <= p2_add_59972_comb;
    p2_add_59973 <= p2_add_59973_comb;
    p2_add_59966 <= p2_add_59966_comb;
    p2_add_59967 <= p2_add_59967_comb;
    p2_add_59968 <= p2_add_59968_comb;
    p2_add_59969 <= p2_add_59969_comb;
    p2_add_59962 <= p2_add_59962_comb;
    p2_add_59963 <= p2_add_59963_comb;
    p2_add_59964 <= p2_add_59964_comb;
    p2_add_59965 <= p2_add_59965_comb;
    p2_add_59958 <= p2_add_59958_comb;
    p2_add_59959 <= p2_add_59959_comb;
    p2_add_59960 <= p2_add_59960_comb;
    p2_add_59961 <= p2_add_59961_comb;
    p2_add_59954 <= p2_add_59954_comb;
    p2_add_59955 <= p2_add_59955_comb;
    p2_add_59956 <= p2_add_59956_comb;
    p2_add_59957 <= p2_add_59957_comb;
    p2_add_59950 <= p2_add_59950_comb;
    p2_add_59951 <= p2_add_59951_comb;
    p2_add_59952 <= p2_add_59952_comb;
    p2_add_59953 <= p2_add_59953_comb;
    p2_add_59946 <= p2_add_59946_comb;
    p2_add_59947 <= p2_add_59947_comb;
    p2_add_59948 <= p2_add_59948_comb;
    p2_add_59949 <= p2_add_59949_comb;
    p2_add_59942 <= p2_add_59942_comb;
    p2_add_59943 <= p2_add_59943_comb;
    p2_add_59944 <= p2_add_59944_comb;
    p2_add_59945 <= p2_add_59945_comb;
    p2_add_59938 <= p2_add_59938_comb;
    p2_add_59939 <= p2_add_59939_comb;
    p2_add_59940 <= p2_add_59940_comb;
    p2_add_59941 <= p2_add_59941_comb;
    p2_add_59934 <= p2_add_59934_comb;
    p2_add_59935 <= p2_add_59935_comb;
    p2_add_59936 <= p2_add_59936_comb;
    p2_add_59937 <= p2_add_59937_comb;
    p2_add_59930 <= p2_add_59930_comb;
    p2_add_59931 <= p2_add_59931_comb;
    p2_add_59932 <= p2_add_59932_comb;
    p2_add_59933 <= p2_add_59933_comb;
    p2_add_59926 <= p2_add_59926_comb;
    p2_add_59927 <= p2_add_59927_comb;
    p2_add_59928 <= p2_add_59928_comb;
    p2_add_59929 <= p2_add_59929_comb;
    p2_add_59922 <= p2_add_59922_comb;
    p2_add_59923 <= p2_add_59923_comb;
    p2_add_59924 <= p2_add_59924_comb;
    p2_add_59925 <= p2_add_59925_comb;
    p2_add_59918 <= p2_add_59918_comb;
    p2_add_59919 <= p2_add_59919_comb;
    p2_add_59920 <= p2_add_59920_comb;
    p2_add_59921 <= p2_add_59921_comb;
    p2_add_59914 <= p2_add_59914_comb;
    p2_add_59915 <= p2_add_59915_comb;
    p2_add_59916 <= p2_add_59916_comb;
    p2_add_59917 <= p2_add_59917_comb;
    p2_add_59910 <= p2_add_59910_comb;
    p2_add_59911 <= p2_add_59911_comb;
    p2_add_59912 <= p2_add_59912_comb;
    p2_add_59913 <= p2_add_59913_comb;
    p2_add_59906 <= p2_add_59906_comb;
    p2_add_59907 <= p2_add_59907_comb;
    p2_add_59908 <= p2_add_59908_comb;
    p2_add_59909 <= p2_add_59909_comb;
    p2_add_59902 <= p2_add_59902_comb;
    p2_add_59903 <= p2_add_59903_comb;
    p2_add_59904 <= p2_add_59904_comb;
    p2_add_59905 <= p2_add_59905_comb;
    p2_add_59898 <= p2_add_59898_comb;
    p2_add_59899 <= p2_add_59899_comb;
    p2_add_59900 <= p2_add_59900_comb;
    p2_add_59901 <= p2_add_59901_comb;
    p2_add_59894 <= p2_add_59894_comb;
    p2_add_59895 <= p2_add_59895_comb;
    p2_add_59896 <= p2_add_59896_comb;
    p2_add_59897 <= p2_add_59897_comb;
    p2_add_59890 <= p2_add_59890_comb;
    p2_add_59891 <= p2_add_59891_comb;
    p2_add_59892 <= p2_add_59892_comb;
    p2_add_59893 <= p2_add_59893_comb;
    p2_add_59886 <= p2_add_59886_comb;
    p2_add_59887 <= p2_add_59887_comb;
    p2_add_59888 <= p2_add_59888_comb;
    p2_add_59889 <= p2_add_59889_comb;
    p2_add_59882 <= p2_add_59882_comb;
    p2_add_59883 <= p2_add_59883_comb;
    p2_add_59884 <= p2_add_59884_comb;
    p2_add_59885 <= p2_add_59885_comb;
    p2_add_59878 <= p2_add_59878_comb;
    p2_add_59879 <= p2_add_59879_comb;
    p2_add_59880 <= p2_add_59880_comb;
    p2_add_59881 <= p2_add_59881_comb;
    p2_add_59874 <= p2_add_59874_comb;
    p2_add_59875 <= p2_add_59875_comb;
    p2_add_59876 <= p2_add_59876_comb;
    p2_add_59877 <= p2_add_59877_comb;
  end

  // ===== Pipe stage 3:
  wire [31:0] p3_add_60646_comb;
  wire [31:0] p3_add_60647_comb;
  wire [31:0] p3_add_60648_comb;
  wire [31:0] p3_add_60649_comb;
  wire [31:0] p3_add_60650_comb;
  wire [31:0] p3_add_60651_comb;
  wire [31:0] p3_add_60652_comb;
  wire [31:0] p3_add_60653_comb;
  wire [31:0] p3_add_60654_comb;
  wire [31:0] p3_add_60655_comb;
  wire [31:0] p3_add_60656_comb;
  wire [31:0] p3_add_60657_comb;
  wire [31:0] p3_add_60658_comb;
  wire [31:0] p3_add_60659_comb;
  wire [31:0] p3_add_60660_comb;
  wire [31:0] p3_add_60661_comb;
  wire [31:0] p3_add_60662_comb;
  wire [31:0] p3_add_60663_comb;
  wire [31:0] p3_add_60664_comb;
  wire [31:0] p3_add_60665_comb;
  wire [31:0] p3_add_60666_comb;
  wire [31:0] p3_add_60667_comb;
  wire [31:0] p3_add_60668_comb;
  wire [31:0] p3_add_60669_comb;
  wire [31:0] p3_add_60670_comb;
  wire [31:0] p3_add_60671_comb;
  wire [31:0] p3_add_60672_comb;
  wire [31:0] p3_add_60673_comb;
  wire [31:0] p3_add_60674_comb;
  wire [31:0] p3_add_60675_comb;
  wire [31:0] p3_add_60676_comb;
  wire [31:0] p3_add_60677_comb;
  wire [31:0] p3_add_60678_comb;
  wire [31:0] p3_add_60679_comb;
  wire [31:0] p3_add_60680_comb;
  wire [31:0] p3_add_60681_comb;
  wire [31:0] p3_add_60682_comb;
  wire [31:0] p3_add_60683_comb;
  wire [31:0] p3_add_60684_comb;
  wire [31:0] p3_add_60685_comb;
  wire [31:0] p3_add_60686_comb;
  wire [31:0] p3_add_60687_comb;
  wire [31:0] p3_add_60688_comb;
  wire [31:0] p3_add_60689_comb;
  wire [31:0] p3_add_60690_comb;
  wire [31:0] p3_add_60691_comb;
  wire [31:0] p3_add_60692_comb;
  wire [31:0] p3_add_60693_comb;
  wire [31:0] p3_add_60694_comb;
  wire [31:0] p3_add_60695_comb;
  wire [31:0] p3_add_60696_comb;
  wire [31:0] p3_add_60697_comb;
  wire [31:0] p3_add_60698_comb;
  wire [31:0] p3_add_60699_comb;
  wire [31:0] p3_add_60700_comb;
  wire [31:0] p3_add_60701_comb;
  wire [31:0] p3_add_60702_comb;
  wire [31:0] p3_add_60703_comb;
  wire [31:0] p3_add_60704_comb;
  wire [31:0] p3_add_60705_comb;
  wire [31:0] p3_add_60706_comb;
  wire [31:0] p3_add_60707_comb;
  wire [31:0] p3_add_60708_comb;
  wire [31:0] p3_add_60709_comb;
  wire [31:0] p3_add_60710_comb;
  wire [31:0] p3_add_60711_comb;
  wire [31:0] p3_add_60712_comb;
  wire [31:0] p3_add_60713_comb;
  wire [31:0] p3_add_60714_comb;
  wire [31:0] p3_add_60715_comb;
  wire [31:0] p3_add_60716_comb;
  wire [31:0] p3_add_60717_comb;
  wire [31:0] p3_add_60718_comb;
  wire [31:0] p3_add_60719_comb;
  wire [31:0] p3_add_60720_comb;
  wire [31:0] p3_add_60721_comb;
  wire [31:0] p3_add_60722_comb;
  wire [31:0] p3_add_60723_comb;
  wire [31:0] p3_add_60724_comb;
  wire [31:0] p3_add_60725_comb;
  wire [31:0] p3_add_60726_comb;
  wire [31:0] p3_add_60727_comb;
  wire [31:0] p3_add_60728_comb;
  wire [31:0] p3_add_60729_comb;
  wire [31:0] p3_add_60730_comb;
  wire [31:0] p3_add_60731_comb;
  wire [31:0] p3_add_60732_comb;
  wire [31:0] p3_add_60733_comb;
  wire [31:0] p3_add_60734_comb;
  wire [31:0] p3_add_60735_comb;
  wire [31:0] p3_add_60736_comb;
  wire [31:0] p3_add_60737_comb;
  wire [31:0] p3_add_60738_comb;
  wire [31:0] p3_add_60739_comb;
  wire [31:0] p3_add_60740_comb;
  wire [31:0] p3_add_60741_comb;
  wire [31:0] p3_add_60742_comb;
  wire [31:0] p3_add_60743_comb;
  wire [31:0] p3_add_60744_comb;
  wire [31:0] p3_add_60745_comb;
  wire [31:0] p3_add_60746_comb;
  wire [31:0] p3_add_60747_comb;
  wire [31:0] p3_add_60748_comb;
  wire [31:0] p3_add_60749_comb;
  wire [31:0] p3_add_60750_comb;
  wire [31:0] p3_add_60751_comb;
  wire [31:0] p3_add_60752_comb;
  wire [31:0] p3_add_60753_comb;
  wire [31:0] p3_add_60754_comb;
  wire [31:0] p3_add_60755_comb;
  wire [31:0] p3_add_60756_comb;
  wire [31:0] p3_add_60757_comb;
  wire [31:0] p3_add_60758_comb;
  wire [31:0] p3_add_60759_comb;
  wire [31:0] p3_add_60760_comb;
  wire [31:0] p3_add_60761_comb;
  wire [31:0] p3_add_60762_comb;
  wire [31:0] p3_add_60763_comb;
  wire [31:0] p3_add_60764_comb;
  wire [31:0] p3_add_60765_comb;
  wire [31:0] p3_add_60766_comb;
  wire [31:0] p3_add_60767_comb;
  wire [31:0] p3_add_60768_comb;
  wire [31:0] p3_add_60769_comb;
  wire [31:0] p3_add_60770_comb;
  wire [31:0] p3_add_60771_comb;
  wire [31:0] p3_add_60772_comb;
  wire [31:0] p3_add_60773_comb;
  wire [31:0] p3_add_60774_comb;
  wire [31:0] p3_add_60775_comb;
  wire [31:0] p3_add_60776_comb;
  wire [31:0] p3_add_60777_comb;
  wire [31:0] p3_add_60778_comb;
  wire [31:0] p3_add_60779_comb;
  wire [31:0] p3_add_60780_comb;
  wire [31:0] p3_add_60781_comb;
  wire [31:0] p3_add_60782_comb;
  wire [31:0] p3_add_60783_comb;
  wire [31:0] p3_add_60784_comb;
  wire [31:0] p3_add_60785_comb;
  wire [31:0] p3_add_60786_comb;
  wire [31:0] p3_add_60787_comb;
  wire [31:0] p3_add_60788_comb;
  wire [31:0] p3_add_60789_comb;
  wire [31:0] p3_add_60790_comb;
  wire [31:0] p3_add_60791_comb;
  wire [31:0] p3_add_60792_comb;
  wire [31:0] p3_add_60793_comb;
  wire [31:0] p3_add_60794_comb;
  wire [31:0] p3_add_60795_comb;
  wire [31:0] p3_add_60796_comb;
  wire [31:0] p3_add_60797_comb;
  wire [31:0] p3_add_60798_comb;
  wire [31:0] p3_add_60799_comb;
  wire [31:0] p3_add_60800_comb;
  wire [31:0] p3_add_60801_comb;
  wire [31:0] p3_add_60802_comb;
  wire [31:0] p3_add_60803_comb;
  wire [31:0] p3_add_60804_comb;
  wire [31:0] p3_add_60805_comb;
  wire [31:0] p3_add_60806_comb;
  wire [31:0] p3_add_60807_comb;
  wire [31:0] p3_add_60808_comb;
  wire [31:0] p3_add_60809_comb;
  wire [31:0] p3_add_60810_comb;
  wire [31:0] p3_add_60811_comb;
  wire [31:0] p3_add_60812_comb;
  wire [31:0] p3_add_60813_comb;
  wire [31:0] p3_add_60814_comb;
  wire [31:0] p3_add_60815_comb;
  wire [31:0] p3_add_60816_comb;
  wire [31:0] p3_add_60817_comb;
  wire [31:0] p3_add_60818_comb;
  wire [31:0] p3_add_60819_comb;
  wire [31:0] p3_add_60820_comb;
  wire [31:0] p3_add_60821_comb;
  wire [31:0] p3_add_60822_comb;
  wire [31:0] p3_add_60823_comb;
  wire [31:0] p3_add_60824_comb;
  wire [31:0] p3_add_60825_comb;
  wire [31:0] p3_add_60826_comb;
  wire [31:0] p3_add_60827_comb;
  wire [31:0] p3_add_60828_comb;
  wire [31:0] p3_add_60829_comb;
  wire [31:0] p3_add_60830_comb;
  wire [31:0] p3_add_60831_comb;
  wire [31:0] p3_add_60832_comb;
  wire [31:0] p3_add_60833_comb;
  wire [31:0] p3_add_60834_comb;
  wire [31:0] p3_add_60835_comb;
  wire [31:0] p3_add_60836_comb;
  wire [31:0] p3_add_60837_comb;
  wire [31:0] p3_array_60838_comb[8];
  wire [31:0] p3_array_60839_comb[8];
  wire [31:0] p3_array_60840_comb[8];
  wire [31:0] p3_array_60841_comb[8];
  wire [31:0] p3_array_60842_comb[8];
  wire [31:0] p3_array_60843_comb[8];
  wire [31:0] p3_array_60844_comb[8];
  wire [31:0] p3_array_60845_comb[8];
  wire [31:0] p3_array_60846_comb[8][8];
  wire [6143:0] p3_tuple_60847_comb;
  assign p3_add_60646_comb = p2_add_59874 + p2_add_59875;
  assign p3_add_60647_comb = p2_add_59876 + p2_add_59877;
  assign p3_add_60648_comb = p2_add_59878 + p2_add_59879;
  assign p3_add_60649_comb = p2_add_59880 + p2_add_59881;
  assign p3_add_60650_comb = p2_add_59882 + p2_add_59883;
  assign p3_add_60651_comb = p2_add_59884 + p2_add_59885;
  assign p3_add_60652_comb = p2_add_59886 + p2_add_59887;
  assign p3_add_60653_comb = p2_add_59888 + p2_add_59889;
  assign p3_add_60654_comb = p2_add_59890 + p2_add_59891;
  assign p3_add_60655_comb = p2_add_59892 + p2_add_59893;
  assign p3_add_60656_comb = p2_add_59894 + p2_add_59895;
  assign p3_add_60657_comb = p2_add_59896 + p2_add_59897;
  assign p3_add_60658_comb = p2_add_59898 + p2_add_59899;
  assign p3_add_60659_comb = p2_add_59900 + p2_add_59901;
  assign p3_add_60660_comb = p2_add_59902 + p2_add_59903;
  assign p3_add_60661_comb = p2_add_59904 + p2_add_59905;
  assign p3_add_60662_comb = p2_add_59906 + p2_add_59907;
  assign p3_add_60663_comb = p2_add_59908 + p2_add_59909;
  assign p3_add_60664_comb = p2_add_59910 + p2_add_59911;
  assign p3_add_60665_comb = p2_add_59912 + p2_add_59913;
  assign p3_add_60666_comb = p2_add_59914 + p2_add_59915;
  assign p3_add_60667_comb = p2_add_59916 + p2_add_59917;
  assign p3_add_60668_comb = p2_add_59918 + p2_add_59919;
  assign p3_add_60669_comb = p2_add_59920 + p2_add_59921;
  assign p3_add_60670_comb = p2_add_59922 + p2_add_59923;
  assign p3_add_60671_comb = p2_add_59924 + p2_add_59925;
  assign p3_add_60672_comb = p2_add_59926 + p2_add_59927;
  assign p3_add_60673_comb = p2_add_59928 + p2_add_59929;
  assign p3_add_60674_comb = p2_add_59930 + p2_add_59931;
  assign p3_add_60675_comb = p2_add_59932 + p2_add_59933;
  assign p3_add_60676_comb = p2_add_59934 + p2_add_59935;
  assign p3_add_60677_comb = p2_add_59936 + p2_add_59937;
  assign p3_add_60678_comb = p2_add_59938 + p2_add_59939;
  assign p3_add_60679_comb = p2_add_59940 + p2_add_59941;
  assign p3_add_60680_comb = p2_add_59942 + p2_add_59943;
  assign p3_add_60681_comb = p2_add_59944 + p2_add_59945;
  assign p3_add_60682_comb = p2_add_59946 + p2_add_59947;
  assign p3_add_60683_comb = p2_add_59948 + p2_add_59949;
  assign p3_add_60684_comb = p2_add_59950 + p2_add_59951;
  assign p3_add_60685_comb = p2_add_59952 + p2_add_59953;
  assign p3_add_60686_comb = p2_add_59954 + p2_add_59955;
  assign p3_add_60687_comb = p2_add_59956 + p2_add_59957;
  assign p3_add_60688_comb = p2_add_59958 + p2_add_59959;
  assign p3_add_60689_comb = p2_add_59960 + p2_add_59961;
  assign p3_add_60690_comb = p2_add_59962 + p2_add_59963;
  assign p3_add_60691_comb = p2_add_59964 + p2_add_59965;
  assign p3_add_60692_comb = p2_add_59966 + p2_add_59967;
  assign p3_add_60693_comb = p2_add_59968 + p2_add_59969;
  assign p3_add_60694_comb = p2_add_59970 + p2_add_59971;
  assign p3_add_60695_comb = p2_add_59972 + p2_add_59973;
  assign p3_add_60696_comb = p2_add_59974 + p2_add_59975;
  assign p3_add_60697_comb = p2_add_59976 + p2_add_59977;
  assign p3_add_60698_comb = p2_add_59978 + p2_add_59979;
  assign p3_add_60699_comb = p2_add_59980 + p2_add_59981;
  assign p3_add_60700_comb = p2_add_59982 + p2_add_59983;
  assign p3_add_60701_comb = p2_add_59984 + p2_add_59985;
  assign p3_add_60702_comb = p2_add_59986 + p2_add_59987;
  assign p3_add_60703_comb = p2_add_59988 + p2_add_59989;
  assign p3_add_60704_comb = p2_add_59990 + p2_add_59991;
  assign p3_add_60705_comb = p2_add_59992 + p2_add_59993;
  assign p3_add_60706_comb = p2_add_59994 + p2_add_59995;
  assign p3_add_60707_comb = p2_add_59996 + p2_add_59997;
  assign p3_add_60708_comb = p2_add_59998 + p2_add_59999;
  assign p3_add_60709_comb = p2_add_60000 + p2_add_60001;
  assign p3_add_60710_comb = p2_add_60002 + p2_add_60003;
  assign p3_add_60711_comb = p2_add_60004 + p2_add_60005;
  assign p3_add_60712_comb = p2_add_60006 + p2_add_60007;
  assign p3_add_60713_comb = p2_add_60008 + p2_add_60009;
  assign p3_add_60714_comb = p2_add_60010 + p2_add_60011;
  assign p3_add_60715_comb = p2_add_60012 + p2_add_60013;
  assign p3_add_60716_comb = p2_add_60014 + p2_add_60015;
  assign p3_add_60717_comb = p2_add_60016 + p2_add_60017;
  assign p3_add_60718_comb = p2_add_60018 + p2_add_60019;
  assign p3_add_60719_comb = p2_add_60020 + p2_add_60021;
  assign p3_add_60720_comb = p2_add_60022 + p2_add_60023;
  assign p3_add_60721_comb = p2_add_60024 + p2_add_60025;
  assign p3_add_60722_comb = p2_add_60026 + p2_add_60027;
  assign p3_add_60723_comb = p2_add_60028 + p2_add_60029;
  assign p3_add_60724_comb = p2_add_60030 + p2_add_60031;
  assign p3_add_60725_comb = p2_add_60032 + p2_add_60033;
  assign p3_add_60726_comb = p2_add_60034 + p2_add_60035;
  assign p3_add_60727_comb = p2_add_60036 + p2_add_60037;
  assign p3_add_60728_comb = p2_add_60038 + p2_add_60039;
  assign p3_add_60729_comb = p2_add_60040 + p2_add_60041;
  assign p3_add_60730_comb = p2_add_60042 + p2_add_60043;
  assign p3_add_60731_comb = p2_add_60044 + p2_add_60045;
  assign p3_add_60732_comb = p2_add_60046 + p2_add_60047;
  assign p3_add_60733_comb = p2_add_60048 + p2_add_60049;
  assign p3_add_60734_comb = p2_add_60050 + p2_add_60051;
  assign p3_add_60735_comb = p2_add_60052 + p2_add_60053;
  assign p3_add_60736_comb = p2_add_60054 + p2_add_60055;
  assign p3_add_60737_comb = p2_add_60056 + p2_add_60057;
  assign p3_add_60738_comb = p2_add_60058 + p2_add_60059;
  assign p3_add_60739_comb = p2_add_60060 + p2_add_60061;
  assign p3_add_60740_comb = p2_add_60062 + p2_add_60063;
  assign p3_add_60741_comb = p2_add_60064 + p2_add_60065;
  assign p3_add_60742_comb = p2_add_60066 + p2_add_60067;
  assign p3_add_60743_comb = p2_add_60068 + p2_add_60069;
  assign p3_add_60744_comb = p2_add_60070 + p2_add_60071;
  assign p3_add_60745_comb = p2_add_60072 + p2_add_60073;
  assign p3_add_60746_comb = p2_add_60074 + p2_add_60075;
  assign p3_add_60747_comb = p2_add_60076 + p2_add_60077;
  assign p3_add_60748_comb = p2_add_60078 + p2_add_60079;
  assign p3_add_60749_comb = p2_add_60080 + p2_add_60081;
  assign p3_add_60750_comb = p2_add_60082 + p2_add_60083;
  assign p3_add_60751_comb = p2_add_60084 + p2_add_60085;
  assign p3_add_60752_comb = p2_add_60086 + p2_add_60087;
  assign p3_add_60753_comb = p2_add_60088 + p2_add_60089;
  assign p3_add_60754_comb = p2_add_60090 + p2_add_60091;
  assign p3_add_60755_comb = p2_add_60092 + p2_add_60093;
  assign p3_add_60756_comb = p2_add_60094 + p2_add_60095;
  assign p3_add_60757_comb = p2_add_60096 + p2_add_60097;
  assign p3_add_60758_comb = p2_add_60098 + p2_add_60099;
  assign p3_add_60759_comb = p2_add_60100 + p2_add_60101;
  assign p3_add_60760_comb = p2_add_60102 + p2_add_60103;
  assign p3_add_60761_comb = p2_add_60104 + p2_add_60105;
  assign p3_add_60762_comb = p2_add_60106 + p2_add_60107;
  assign p3_add_60763_comb = p2_add_60108 + p2_add_60109;
  assign p3_add_60764_comb = p2_add_60110 + p2_add_60111;
  assign p3_add_60765_comb = p2_add_60112 + p2_add_60113;
  assign p3_add_60766_comb = p2_add_60114 + p2_add_60115;
  assign p3_add_60767_comb = p2_add_60116 + p2_add_60117;
  assign p3_add_60768_comb = p2_add_60118 + p2_add_60119;
  assign p3_add_60769_comb = p2_add_60120 + p2_add_60121;
  assign p3_add_60770_comb = p2_add_60122 + p2_add_60123;
  assign p3_add_60771_comb = p2_add_60124 + p2_add_60125;
  assign p3_add_60772_comb = p2_add_60126 + p2_add_60127;
  assign p3_add_60773_comb = p2_add_60128 + p2_add_60129;
  assign p3_add_60774_comb = p3_add_60646_comb + p3_add_60647_comb;
  assign p3_add_60775_comb = p3_add_60648_comb + p3_add_60649_comb;
  assign p3_add_60776_comb = p3_add_60650_comb + p3_add_60651_comb;
  assign p3_add_60777_comb = p3_add_60652_comb + p3_add_60653_comb;
  assign p3_add_60778_comb = p3_add_60654_comb + p3_add_60655_comb;
  assign p3_add_60779_comb = p3_add_60656_comb + p3_add_60657_comb;
  assign p3_add_60780_comb = p3_add_60658_comb + p3_add_60659_comb;
  assign p3_add_60781_comb = p3_add_60660_comb + p3_add_60661_comb;
  assign p3_add_60782_comb = p3_add_60662_comb + p3_add_60663_comb;
  assign p3_add_60783_comb = p3_add_60664_comb + p3_add_60665_comb;
  assign p3_add_60784_comb = p3_add_60666_comb + p3_add_60667_comb;
  assign p3_add_60785_comb = p3_add_60668_comb + p3_add_60669_comb;
  assign p3_add_60786_comb = p3_add_60670_comb + p3_add_60671_comb;
  assign p3_add_60787_comb = p3_add_60672_comb + p3_add_60673_comb;
  assign p3_add_60788_comb = p3_add_60674_comb + p3_add_60675_comb;
  assign p3_add_60789_comb = p3_add_60676_comb + p3_add_60677_comb;
  assign p3_add_60790_comb = p3_add_60678_comb + p3_add_60679_comb;
  assign p3_add_60791_comb = p3_add_60680_comb + p3_add_60681_comb;
  assign p3_add_60792_comb = p3_add_60682_comb + p3_add_60683_comb;
  assign p3_add_60793_comb = p3_add_60684_comb + p3_add_60685_comb;
  assign p3_add_60794_comb = p3_add_60686_comb + p3_add_60687_comb;
  assign p3_add_60795_comb = p3_add_60688_comb + p3_add_60689_comb;
  assign p3_add_60796_comb = p3_add_60690_comb + p3_add_60691_comb;
  assign p3_add_60797_comb = p3_add_60692_comb + p3_add_60693_comb;
  assign p3_add_60798_comb = p3_add_60694_comb + p3_add_60695_comb;
  assign p3_add_60799_comb = p3_add_60696_comb + p3_add_60697_comb;
  assign p3_add_60800_comb = p3_add_60698_comb + p3_add_60699_comb;
  assign p3_add_60801_comb = p3_add_60700_comb + p3_add_60701_comb;
  assign p3_add_60802_comb = p3_add_60702_comb + p3_add_60703_comb;
  assign p3_add_60803_comb = p3_add_60704_comb + p3_add_60705_comb;
  assign p3_add_60804_comb = p3_add_60706_comb + p3_add_60707_comb;
  assign p3_add_60805_comb = p3_add_60708_comb + p3_add_60709_comb;
  assign p3_add_60806_comb = p3_add_60710_comb + p3_add_60711_comb;
  assign p3_add_60807_comb = p3_add_60712_comb + p3_add_60713_comb;
  assign p3_add_60808_comb = p3_add_60714_comb + p3_add_60715_comb;
  assign p3_add_60809_comb = p3_add_60716_comb + p3_add_60717_comb;
  assign p3_add_60810_comb = p3_add_60718_comb + p3_add_60719_comb;
  assign p3_add_60811_comb = p3_add_60720_comb + p3_add_60721_comb;
  assign p3_add_60812_comb = p3_add_60722_comb + p3_add_60723_comb;
  assign p3_add_60813_comb = p3_add_60724_comb + p3_add_60725_comb;
  assign p3_add_60814_comb = p3_add_60726_comb + p3_add_60727_comb;
  assign p3_add_60815_comb = p3_add_60728_comb + p3_add_60729_comb;
  assign p3_add_60816_comb = p3_add_60730_comb + p3_add_60731_comb;
  assign p3_add_60817_comb = p3_add_60732_comb + p3_add_60733_comb;
  assign p3_add_60818_comb = p3_add_60734_comb + p3_add_60735_comb;
  assign p3_add_60819_comb = p3_add_60736_comb + p3_add_60737_comb;
  assign p3_add_60820_comb = p3_add_60738_comb + p3_add_60739_comb;
  assign p3_add_60821_comb = p3_add_60740_comb + p3_add_60741_comb;
  assign p3_add_60822_comb = p3_add_60742_comb + p3_add_60743_comb;
  assign p3_add_60823_comb = p3_add_60744_comb + p3_add_60745_comb;
  assign p3_add_60824_comb = p3_add_60746_comb + p3_add_60747_comb;
  assign p3_add_60825_comb = p3_add_60748_comb + p3_add_60749_comb;
  assign p3_add_60826_comb = p3_add_60750_comb + p3_add_60751_comb;
  assign p3_add_60827_comb = p3_add_60752_comb + p3_add_60753_comb;
  assign p3_add_60828_comb = p3_add_60754_comb + p3_add_60755_comb;
  assign p3_add_60829_comb = p3_add_60756_comb + p3_add_60757_comb;
  assign p3_add_60830_comb = p3_add_60758_comb + p3_add_60759_comb;
  assign p3_add_60831_comb = p3_add_60760_comb + p3_add_60761_comb;
  assign p3_add_60832_comb = p3_add_60762_comb + p3_add_60763_comb;
  assign p3_add_60833_comb = p3_add_60764_comb + p3_add_60765_comb;
  assign p3_add_60834_comb = p3_add_60766_comb + p3_add_60767_comb;
  assign p3_add_60835_comb = p3_add_60768_comb + p3_add_60769_comb;
  assign p3_add_60836_comb = p3_add_60770_comb + p3_add_60771_comb;
  assign p3_add_60837_comb = p3_add_60772_comb + p3_add_60773_comb;
  assign p3_array_60838_comb[0] = p3_add_60774_comb;
  assign p3_array_60838_comb[1] = p3_add_60775_comb;
  assign p3_array_60838_comb[2] = p3_add_60776_comb;
  assign p3_array_60838_comb[3] = p3_add_60777_comb;
  assign p3_array_60838_comb[4] = p3_add_60778_comb;
  assign p3_array_60838_comb[5] = p3_add_60779_comb;
  assign p3_array_60838_comb[6] = p3_add_60780_comb;
  assign p3_array_60838_comb[7] = p3_add_60781_comb;
  assign p3_array_60839_comb[0] = p3_add_60782_comb;
  assign p3_array_60839_comb[1] = p3_add_60783_comb;
  assign p3_array_60839_comb[2] = p3_add_60784_comb;
  assign p3_array_60839_comb[3] = p3_add_60785_comb;
  assign p3_array_60839_comb[4] = p3_add_60786_comb;
  assign p3_array_60839_comb[5] = p3_add_60787_comb;
  assign p3_array_60839_comb[6] = p3_add_60788_comb;
  assign p3_array_60839_comb[7] = p3_add_60789_comb;
  assign p3_array_60840_comb[0] = p3_add_60790_comb;
  assign p3_array_60840_comb[1] = p3_add_60791_comb;
  assign p3_array_60840_comb[2] = p3_add_60792_comb;
  assign p3_array_60840_comb[3] = p3_add_60793_comb;
  assign p3_array_60840_comb[4] = p3_add_60794_comb;
  assign p3_array_60840_comb[5] = p3_add_60795_comb;
  assign p3_array_60840_comb[6] = p3_add_60796_comb;
  assign p3_array_60840_comb[7] = p3_add_60797_comb;
  assign p3_array_60841_comb[0] = p3_add_60798_comb;
  assign p3_array_60841_comb[1] = p3_add_60799_comb;
  assign p3_array_60841_comb[2] = p3_add_60800_comb;
  assign p3_array_60841_comb[3] = p3_add_60801_comb;
  assign p3_array_60841_comb[4] = p3_add_60802_comb;
  assign p3_array_60841_comb[5] = p3_add_60803_comb;
  assign p3_array_60841_comb[6] = p3_add_60804_comb;
  assign p3_array_60841_comb[7] = p3_add_60805_comb;
  assign p3_array_60842_comb[0] = p3_add_60806_comb;
  assign p3_array_60842_comb[1] = p3_add_60807_comb;
  assign p3_array_60842_comb[2] = p3_add_60808_comb;
  assign p3_array_60842_comb[3] = p3_add_60809_comb;
  assign p3_array_60842_comb[4] = p3_add_60810_comb;
  assign p3_array_60842_comb[5] = p3_add_60811_comb;
  assign p3_array_60842_comb[6] = p3_add_60812_comb;
  assign p3_array_60842_comb[7] = p3_add_60813_comb;
  assign p3_array_60843_comb[0] = p3_add_60814_comb;
  assign p3_array_60843_comb[1] = p3_add_60815_comb;
  assign p3_array_60843_comb[2] = p3_add_60816_comb;
  assign p3_array_60843_comb[3] = p3_add_60817_comb;
  assign p3_array_60843_comb[4] = p3_add_60818_comb;
  assign p3_array_60843_comb[5] = p3_add_60819_comb;
  assign p3_array_60843_comb[6] = p3_add_60820_comb;
  assign p3_array_60843_comb[7] = p3_add_60821_comb;
  assign p3_array_60844_comb[0] = p3_add_60822_comb;
  assign p3_array_60844_comb[1] = p3_add_60823_comb;
  assign p3_array_60844_comb[2] = p3_add_60824_comb;
  assign p3_array_60844_comb[3] = p3_add_60825_comb;
  assign p3_array_60844_comb[4] = p3_add_60826_comb;
  assign p3_array_60844_comb[5] = p3_add_60827_comb;
  assign p3_array_60844_comb[6] = p3_add_60828_comb;
  assign p3_array_60844_comb[7] = p3_add_60829_comb;
  assign p3_array_60845_comb[0] = p3_add_60830_comb;
  assign p3_array_60845_comb[1] = p3_add_60831_comb;
  assign p3_array_60845_comb[2] = p3_add_60832_comb;
  assign p3_array_60845_comb[3] = p3_add_60833_comb;
  assign p3_array_60845_comb[4] = p3_add_60834_comb;
  assign p3_array_60845_comb[5] = p3_add_60835_comb;
  assign p3_array_60845_comb[6] = p3_add_60836_comb;
  assign p3_array_60845_comb[7] = p3_add_60837_comb;
  assign p3_array_60846_comb[0] = p3_array_60838_comb;
  assign p3_array_60846_comb[1] = p3_array_60839_comb;
  assign p3_array_60846_comb[2] = p3_array_60840_comb;
  assign p3_array_60846_comb[3] = p3_array_60841_comb;
  assign p3_array_60846_comb[4] = p3_array_60842_comb;
  assign p3_array_60846_comb[5] = p3_array_60843_comb;
  assign p3_array_60846_comb[6] = p3_array_60844_comb;
  assign p3_array_60846_comb[7] = p3_array_60845_comb;
  assign p3_tuple_60847_comb = {{{p2_a[7][7], p2_a[7][6], p2_a[7][5], p2_a[7][4], p2_a[7][3], p2_a[7][2], p2_a[7][1], p2_a[7][0]}, {p2_a[6][7], p2_a[6][6], p2_a[6][5], p2_a[6][4], p2_a[6][3], p2_a[6][2], p2_a[6][1], p2_a[6][0]}, {p2_a[5][7], p2_a[5][6], p2_a[5][5], p2_a[5][4], p2_a[5][3], p2_a[5][2], p2_a[5][1], p2_a[5][0]}, {p2_a[4][7], p2_a[4][6], p2_a[4][5], p2_a[4][4], p2_a[4][3], p2_a[4][2], p2_a[4][1], p2_a[4][0]}, {p2_a[3][7], p2_a[3][6], p2_a[3][5], p2_a[3][4], p2_a[3][3], p2_a[3][2], p2_a[3][1], p2_a[3][0]}, {p2_a[2][7], p2_a[2][6], p2_a[2][5], p2_a[2][4], p2_a[2][3], p2_a[2][2], p2_a[2][1], p2_a[2][0]}, {p2_a[1][7], p2_a[1][6], p2_a[1][5], p2_a[1][4], p2_a[1][3], p2_a[1][2], p2_a[1][1], p2_a[1][0]}, {p2_a[0][7], p2_a[0][6], p2_a[0][5], p2_a[0][4], p2_a[0][3], p2_a[0][2], p2_a[0][1], p2_a[0][0]}}, {{p2_b[7][7], p2_b[7][6], p2_b[7][5], p2_b[7][4], p2_b[7][3], p2_b[7][2], p2_b[7][1], p2_b[7][0]}, {p2_b[6][7], p2_b[6][6], p2_b[6][5], p2_b[6][4], p2_b[6][3], p2_b[6][2], p2_b[6][1], p2_b[6][0]}, {p2_b[5][7], p2_b[5][6], p2_b[5][5], p2_b[5][4], p2_b[5][3], p2_b[5][2], p2_b[5][1], p2_b[5][0]}, {p2_b[4][7], p2_b[4][6], p2_b[4][5], p2_b[4][4], p2_b[4][3], p2_b[4][2], p2_b[4][1], p2_b[4][0]}, {p2_b[3][7], p2_b[3][6], p2_b[3][5], p2_b[3][4], p2_b[3][3], p2_b[3][2], p2_b[3][1], p2_b[3][0]}, {p2_b[2][7], p2_b[2][6], p2_b[2][5], p2_b[2][4], p2_b[2][3], p2_b[2][2], p2_b[2][1], p2_b[2][0]}, {p2_b[1][7], p2_b[1][6], p2_b[1][5], p2_b[1][4], p2_b[1][3], p2_b[1][2], p2_b[1][1], p2_b[1][0]}, {p2_b[0][7], p2_b[0][6], p2_b[0][5], p2_b[0][4], p2_b[0][3], p2_b[0][2], p2_b[0][1], p2_b[0][0]}}, {{p3_array_60846_comb[7][7], p3_array_60846_comb[7][6], p3_array_60846_comb[7][5], p3_array_60846_comb[7][4], p3_array_60846_comb[7][3], p3_array_60846_comb[7][2], p3_array_60846_comb[7][1], p3_array_60846_comb[7][0]}, {p3_array_60846_comb[6][7], p3_array_60846_comb[6][6], p3_array_60846_comb[6][5], p3_array_60846_comb[6][4], p3_array_60846_comb[6][3], p3_array_60846_comb[6][2], p3_array_60846_comb[6][1], p3_array_60846_comb[6][0]}, {p3_array_60846_comb[5][7], p3_array_60846_comb[5][6], p3_array_60846_comb[5][5], p3_array_60846_comb[5][4], p3_array_60846_comb[5][3], p3_array_60846_comb[5][2], p3_array_60846_comb[5][1], p3_array_60846_comb[5][0]}, {p3_array_60846_comb[4][7], p3_array_60846_comb[4][6], p3_array_60846_comb[4][5], p3_array_60846_comb[4][4], p3_array_60846_comb[4][3], p3_array_60846_comb[4][2], p3_array_60846_comb[4][1], p3_array_60846_comb[4][0]}, {p3_array_60846_comb[3][7], p3_array_60846_comb[3][6], p3_array_60846_comb[3][5], p3_array_60846_comb[3][4], p3_array_60846_comb[3][3], p3_array_60846_comb[3][2], p3_array_60846_comb[3][1], p3_array_60846_comb[3][0]}, {p3_array_60846_comb[2][7], p3_array_60846_comb[2][6], p3_array_60846_comb[2][5], p3_array_60846_comb[2][4], p3_array_60846_comb[2][3], p3_array_60846_comb[2][2], p3_array_60846_comb[2][1], p3_array_60846_comb[2][0]}, {p3_array_60846_comb[1][7], p3_array_60846_comb[1][6], p3_array_60846_comb[1][5], p3_array_60846_comb[1][4], p3_array_60846_comb[1][3], p3_array_60846_comb[1][2], p3_array_60846_comb[1][1], p3_array_60846_comb[1][0]}, {p3_array_60846_comb[0][7], p3_array_60846_comb[0][6], p3_array_60846_comb[0][5], p3_array_60846_comb[0][4], p3_array_60846_comb[0][3], p3_array_60846_comb[0][2], p3_array_60846_comb[0][1], p3_array_60846_comb[0][0]}}};

  // Registers for pipe stage 3:
  reg [6143:0] p3_tuple_60847;
  always_ff @ (posedge clk) begin
    p3_tuple_60847 <= p3_tuple_60847_comb;
  end
  assign out = p3_tuple_60847;
endmodule
