module xls_test(
  input wire clk,
  input wire [511:0] message,
  output wire [255:0] out
);
  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [511:0] p0_message;
  always_ff @ (posedge clk) begin
    p0_message <= message;
  end

  // ===== Pipe stage 1:
  wire [28:0] p1_add_62796_comb;
  wire [30:0] p1_add_62800_comb;
  wire [29:0] p1_add_62803_comb;
  assign p1_add_62796_comb = p0_message[511:483] + 29'h1e6e_fdad;
  assign p1_add_62800_comb = {p1_add_62796_comb, p0_message[482:481]} + 31'h52a7_fa9d;
  assign p1_add_62803_comb = p0_message[479:450] + 30'h242e_c78f;

  // Registers for pipe stage 1:
  reg [511:0] p1_message;
  reg [28:0] p1_add_62796;
  reg [30:0] p1_add_62800;
  reg [29:0] p1_add_62803;
  always_ff @ (posedge clk) begin
    p1_message <= p0_message;
    p1_add_62796 <= p1_add_62796_comb;
    p1_add_62800 <= p1_add_62800_comb;
    p1_add_62803 <= p1_add_62803_comb;
  end

  // ===== Pipe stage 2:
  wire p2_bit_slice_62812_comb;
  wire [31:0] p2_concat_62813_comb;
  wire [31:0] p2_add_62840_comb;
  wire [31:0] p2_add_62842_comb;
  wire [30:0] p2_add_62845_comb;
  assign p2_bit_slice_62812_comb = p1_message[480];
  assign p2_concat_62813_comb = {p1_add_62800, p2_bit_slice_62812_comb};
  assign p2_add_62840_comb = (p2_concat_62813_comb & 32'h510e_527f ^ ~(p2_concat_62813_comb | 32'h64fa_9773)) + {p1_add_62803, p1_message[449:448]};
  assign p2_add_62842_comb = p2_add_62840_comb + {{p1_add_62800[4:0], p2_bit_slice_62812_comb} ^ p1_add_62800[9:4] ^ p1_add_62800[23:18], p1_add_62800[30:26] ^ {p1_add_62800[3:0], p2_bit_slice_62812_comb} ^ p1_add_62800[17:13], p1_add_62800[25:12] ^ p1_add_62800[30:17] ^ {p1_add_62800[12:0], p2_bit_slice_62812_comb}, p1_add_62800[11:5] ^ p1_add_62800[16:10] ^ p1_add_62800[30:24]};
  assign p2_add_62845_comb = p2_add_62842_comb[31:1] + 31'h1e37_79b9;

  // Registers for pipe stage 2:
  reg [511:0] p2_message;
  reg p2_bit_slice_62812;
  reg [31:0] p2_concat_62813;
  reg [31:0] p2_add_62842;
  reg [28:0] p2_add_62796;
  reg [30:0] p2_add_62800;
  reg [30:0] p2_add_62845;
  always_ff @ (posedge clk) begin
    p2_message <= p1_message;
    p2_bit_slice_62812 <= p2_bit_slice_62812_comb;
    p2_concat_62813 <= p2_concat_62813_comb;
    p2_add_62842 <= p2_add_62842_comb;
    p2_add_62796 <= p1_add_62796;
    p2_add_62800 <= p1_add_62800;
    p2_add_62845 <= p2_add_62845_comb;
  end

  // ===== Pipe stage 3:
  wire [31:0] p3_concat_62866_comb;
  wire [31:0] p3_bit_slice_62886_comb;
  wire [31:0] p3_add_62908_comb;
  wire [31:0] p3_add_62890_comb;
  wire [31:0] p3_add_62891_comb;
  wire [31:0] p3_and_62911_comb;
  wire [31:0] p3_add_62892_comb;
  wire [31:0] p3_add_62896_comb;
  wire [31:0] p3_add_62931_comb;
  wire [31:0] p3_nor_62900_comb;
  wire [31:0] p3_concat_62904_comb;
  wire [31:0] p3_add_62933_comb;
  wire [29:0] p3_add_62901_comb;
  assign p3_concat_62866_comb = {p2_add_62845, p2_add_62842[0]};
  assign p3_bit_slice_62886_comb = p2_message[447:416];
  assign p3_add_62908_comb = {p2_add_62796, p2_message[482:480]} + 32'h0890_9ae5;
  assign p3_add_62890_comb = p3_bit_slice_62886_comb + ({p2_add_62845 & p2_add_62800, p2_add_62842[0] & p2_bit_slice_62812} ^ ~(p3_concat_62866_comb | 32'haef1_ad80));
  assign p3_add_62891_comb = {{p2_add_62845[4:0], p2_add_62842[0]} ^ p2_add_62845[9:4] ^ p2_add_62845[23:18], p2_add_62845[30:26] ^ {p2_add_62845[3:0], p2_add_62842[0]} ^ p2_add_62845[17:13], p2_add_62845[25:12] ^ p2_add_62845[30:17] ^ {p2_add_62845[12:0], p2_add_62842[0]}, p2_add_62845[11:5] ^ p2_add_62845[16:10] ^ p2_add_62845[30:24]} + 32'h50c6_645b;
  assign p3_and_62911_comb = p3_add_62908_comb & 32'h6a09_e667;
  assign p3_add_62892_comb = p3_add_62890_comb + p3_add_62891_comb;
  assign p3_add_62896_comb = p3_add_62892_comb + 32'hbb67_ae85;
  assign p3_add_62931_comb = (p3_and_62911_comb ^ p3_add_62908_comb & 32'hbb67_ae85 ^ 32'h2a01_a605) + p2_add_62842;
  assign p3_nor_62900_comb = ~(p3_add_62896_comb | {~p2_add_62800, ~p2_bit_slice_62812});
  assign p3_concat_62904_comb = {~p2_add_62845, ~p2_add_62842[0]};
  assign p3_add_62933_comb = p3_add_62931_comb + {p3_add_62908_comb[1:0] ^ p3_add_62908_comb[12:11] ^ p3_add_62908_comb[21:20], p3_add_62908_comb[31:21] ^ p3_add_62908_comb[10:0] ^ p3_add_62908_comb[19:9], p3_add_62908_comb[20:12] ^ p3_add_62908_comb[31:23] ^ p3_add_62908_comb[8:0], p3_add_62908_comb[11:2] ^ p3_add_62908_comb[22:13] ^ p3_add_62908_comb[31:22]};
  assign p3_add_62901_comb = p2_message[415:386] + 30'h0eb1_0b89;

  // Registers for pipe stage 3:
  reg [511:0] p3_message;
  reg [31:0] p3_concat_62813;
  reg [31:0] p3_concat_62866;
  reg [31:0] p3_bit_slice_62886;
  reg [31:0] p3_add_62892;
  reg [31:0] p3_nor_62900;
  reg [31:0] p3_concat_62904;
  reg [31:0] p3_and_62911;
  reg [31:0] p3_add_62933;
  reg [31:0] p3_add_62896;
  reg [29:0] p3_add_62901;
  reg [31:0] p3_add_62908;
  always_ff @ (posedge clk) begin
    p3_message <= p2_message;
    p3_concat_62813 <= p2_concat_62813;
    p3_concat_62866 <= p3_concat_62866_comb;
    p3_bit_slice_62886 <= p3_bit_slice_62886_comb;
    p3_add_62892 <= p3_add_62892_comb;
    p3_nor_62900 <= p3_nor_62900_comb;
    p3_concat_62904 <= p3_concat_62904_comb;
    p3_and_62911 <= p3_and_62911_comb;
    p3_add_62933 <= p3_add_62933_comb;
    p3_add_62896 <= p3_add_62896_comb;
    p3_add_62901 <= p3_add_62901_comb;
    p3_add_62908 <= p3_add_62908_comb;
  end

  // ===== Pipe stage 4:
  wire [31:0] p4_add_62978_comb;
  wire [31:0] p4_and_62989_comb;
  wire [31:0] p4_add_62980_comb;
  wire [31:0] p4_bit_slice_62984_comb;
  wire [31:0] p4_add_62982_comb;
  wire [31:0] p4_add_62986_comb;
  wire [31:0] p4_add_63008_comb;
  wire [31:0] p4_nor_62983_comb;
  wire [31:0] p4_add_62987_comb;
  wire [31:0] p4_add_63010_comb;
  assign p4_add_62978_comb = (p3_add_62896 & p3_concat_62866 ^ p3_nor_62900) + {p3_add_62901, p3_message[385:384]};
  assign p4_and_62989_comb = p3_add_62933 & p3_add_62908;
  assign p4_add_62980_comb = p4_add_62978_comb + {p3_add_62896[5:0] ^ p3_add_62896[10:5] ^ p3_add_62896[24:19], p3_add_62896[31:27] ^ p3_add_62896[4:0] ^ p3_add_62896[18:14], p3_add_62896[26:13] ^ p3_add_62896[31:18] ^ p3_add_62896[13:0], p3_add_62896[12:6] ^ p3_add_62896[17:11] ^ p3_add_62896[31:25]};
  assign p4_bit_slice_62984_comb = p3_message[383:352];
  assign p4_add_62982_comb = p4_add_62980_comb + 32'h6a09_e667;
  assign p4_add_62986_comb = p4_bit_slice_62984_comb + 32'h3956_c25b;
  assign p4_add_63008_comb = (p4_and_62989_comb ^ p3_add_62933 & 32'h6a09_e667 ^ p3_and_62911) + p3_add_62892;
  assign p4_nor_62983_comb = ~(p4_add_62982_comb | p3_concat_62904);
  assign p4_add_62987_comb = p3_concat_62813 + p4_add_62986_comb;
  assign p4_add_63010_comb = p4_add_63008_comb + {p3_add_62933[1:0] ^ p3_add_62933[12:11] ^ p3_add_62933[21:20], p3_add_62933[31:21] ^ p3_add_62933[10:0] ^ p3_add_62933[19:9], p3_add_62933[20:12] ^ p3_add_62933[31:23] ^ p3_add_62933[8:0], p3_add_62933[11:2] ^ p3_add_62933[22:13] ^ p3_add_62933[31:22]};

  // Registers for pipe stage 4:
  reg [511:0] p4_message;
  reg [31:0] p4_concat_62866;
  reg [31:0] p4_bit_slice_62886;
  reg [31:0] p4_add_62980;
  reg [31:0] p4_nor_62983;
  reg [31:0] p4_bit_slice_62984;
  reg [31:0] p4_add_62987;
  reg [31:0] p4_add_62933;
  reg [31:0] p4_and_62989;
  reg [31:0] p4_add_63010;
  reg [31:0] p4_add_62896;
  reg [31:0] p4_add_62982;
  reg [31:0] p4_add_62908;
  always_ff @ (posedge clk) begin
    p4_message <= p3_message;
    p4_concat_62866 <= p3_concat_62866;
    p4_bit_slice_62886 <= p3_bit_slice_62886;
    p4_add_62980 <= p4_add_62980_comb;
    p4_nor_62983 <= p4_nor_62983_comb;
    p4_bit_slice_62984 <= p4_bit_slice_62984_comb;
    p4_add_62987 <= p4_add_62987_comb;
    p4_add_62933 <= p3_add_62933;
    p4_and_62989 <= p4_and_62989_comb;
    p4_add_63010 <= p4_add_63010_comb;
    p4_add_62896 <= p3_add_62896;
    p4_add_62982 <= p4_add_62982_comb;
    p4_add_62908 <= p3_add_62908;
  end

  // ===== Pipe stage 5:
  wire [31:0] p5_and_63063_comb;
  wire [31:0] p5_add_63056_comb;
  wire [31:0] p5_bit_slice_63059_comb;
  wire [31:0] p5_add_63057_comb;
  wire [31:0] p5_add_63061_comb;
  wire [31:0] p5_add_63082_comb;
  wire [31:0] p5_add_63058_comb;
  wire [31:0] p5_add_63062_comb;
  wire [31:0] p5_add_63084_comb;
  assign p5_and_63063_comb = p4_add_63010 & p4_add_62933;
  assign p5_add_63056_comb = {p4_add_62982[5:0] ^ p4_add_62982[10:5] ^ p4_add_62982[24:19], p4_add_62982[31:27] ^ p4_add_62982[4:0] ^ p4_add_62982[18:14], p4_add_62982[26:13] ^ p4_add_62982[31:18] ^ p4_add_62982[13:0], p4_add_62982[12:6] ^ p4_add_62982[17:11] ^ p4_add_62982[31:25]} + (p4_add_62982 & p4_add_62896 ^ p4_nor_62983);
  assign p5_bit_slice_63059_comb = p4_message[351:320];
  assign p5_add_63057_comb = p5_add_63056_comb + p4_add_62987;
  assign p5_add_63061_comb = p5_bit_slice_63059_comb + 32'h59f1_11f1;
  assign p5_add_63082_comb = (p5_and_63063_comb ^ p4_add_63010 & p4_add_62908 ^ p4_and_62989) + p4_add_62980;
  assign p5_add_63058_comb = p5_add_63057_comb + p4_add_62908;
  assign p5_add_63062_comb = p4_concat_62866 + p5_add_63061_comb;
  assign p5_add_63084_comb = p5_add_63082_comb + {p4_add_63010[1:0] ^ p4_add_63010[12:11] ^ p4_add_63010[21:20], p4_add_63010[31:21] ^ p4_add_63010[10:0] ^ p4_add_63010[19:9], p4_add_63010[20:12] ^ p4_add_63010[31:23] ^ p4_add_63010[8:0], p4_add_63010[11:2] ^ p4_add_63010[22:13] ^ p4_add_63010[31:22]};

  // Registers for pipe stage 5:
  reg [511:0] p5_message;
  reg [31:0] p5_bit_slice_62886;
  reg [31:0] p5_bit_slice_62984;
  reg [31:0] p5_add_63057;
  reg [31:0] p5_add_63058;
  reg [31:0] p5_bit_slice_63059;
  reg [31:0] p5_add_63062;
  reg [31:0] p5_add_62933;
  reg [31:0] p5_add_63010;
  reg [31:0] p5_and_63063;
  reg [31:0] p5_add_63084;
  reg [31:0] p5_add_62896;
  reg [31:0] p5_add_62982;
  always_ff @ (posedge clk) begin
    p5_message <= p4_message;
    p5_bit_slice_62886 <= p4_bit_slice_62886;
    p5_bit_slice_62984 <= p4_bit_slice_62984;
    p5_add_63057 <= p5_add_63057_comb;
    p5_add_63058 <= p5_add_63058_comb;
    p5_bit_slice_63059 <= p5_bit_slice_63059_comb;
    p5_add_63062 <= p5_add_63062_comb;
    p5_add_62933 <= p4_add_62933;
    p5_add_63010 <= p4_add_63010;
    p5_and_63063 <= p5_and_63063_comb;
    p5_add_63084 <= p5_add_63084_comb;
    p5_add_62896 <= p4_add_62896;
    p5_add_62982 <= p4_add_62982;
  end

  // ===== Pipe stage 6:
  wire [31:0] p6_and_63141_comb;
  wire [31:0] p6_add_63132_comb;
  wire [29:0] p6_add_63137_comb;
  wire [31:0] p6_add_63133_comb;
  wire [31:0] p6_add_63160_comb;
  wire [31:0] p6_add_63134_comb;
  wire [31:0] p6_add_63140_comb;
  wire [31:0] p6_add_63162_comb;
  assign p6_and_63141_comb = p5_add_63084 & p5_add_63010;
  assign p6_add_63132_comb = {p5_add_63058[5:0] ^ p5_add_63058[10:5] ^ p5_add_63058[24:19], p5_add_63058[31:27] ^ p5_add_63058[4:0] ^ p5_add_63058[18:14], p5_add_63058[26:13] ^ p5_add_63058[31:18] ^ p5_add_63058[13:0], p5_add_63058[12:6] ^ p5_add_63058[17:11] ^ p5_add_63058[31:25]} + (p5_add_63058 & p5_add_62982 ^ ~(p5_add_63058 | ~p5_add_62896));
  assign p6_add_63137_comb = p5_message[319:290] + 30'h248f_e0a9;
  assign p6_add_63133_comb = p6_add_63132_comb + p5_add_63062;
  assign p6_add_63160_comb = (p6_and_63141_comb ^ p5_add_63084 & p5_add_62933 ^ p5_and_63063) + p5_add_63057;
  assign p6_add_63134_comb = p6_add_63133_comb + p5_add_62933;
  assign p6_add_63140_comb = {p6_add_63137_comb, p5_message[289:288]} + p5_add_62896;
  assign p6_add_63162_comb = p6_add_63160_comb + {p5_add_63084[1:0] ^ p5_add_63084[12:11] ^ p5_add_63084[21:20], p5_add_63084[31:21] ^ p5_add_63084[10:0] ^ p5_add_63084[19:9], p5_add_63084[20:12] ^ p5_add_63084[31:23] ^ p5_add_63084[8:0], p5_add_63084[11:2] ^ p5_add_63084[22:13] ^ p5_add_63084[31:22]};

  // Registers for pipe stage 6:
  reg [511:0] p6_message;
  reg [31:0] p6_bit_slice_62886;
  reg [31:0] p6_bit_slice_62984;
  reg [31:0] p6_add_63058;
  reg [31:0] p6_bit_slice_63059;
  reg [31:0] p6_add_63133;
  reg [31:0] p6_add_63134;
  reg [31:0] p6_add_63140;
  reg [31:0] p6_add_63010;
  reg [31:0] p6_add_63084;
  reg [31:0] p6_and_63141;
  reg [31:0] p6_add_63162;
  reg [31:0] p6_add_62982;
  always_ff @ (posedge clk) begin
    p6_message <= p5_message;
    p6_bit_slice_62886 <= p5_bit_slice_62886;
    p6_bit_slice_62984 <= p5_bit_slice_62984;
    p6_add_63058 <= p5_add_63058;
    p6_bit_slice_63059 <= p5_bit_slice_63059;
    p6_add_63133 <= p6_add_63133_comb;
    p6_add_63134 <= p6_add_63134_comb;
    p6_add_63140 <= p6_add_63140_comb;
    p6_add_63010 <= p5_add_63010;
    p6_add_63084 <= p5_add_63084;
    p6_and_63141 <= p6_and_63141_comb;
    p6_add_63162 <= p6_add_63162_comb;
    p6_add_62982 <= p5_add_62982;
  end

  // ===== Pipe stage 7:
  wire [31:0] p7_and_63217_comb;
  wire [31:0] p7_add_63210_comb;
  wire [31:0] p7_bit_slice_63213_comb;
  wire [31:0] p7_add_63211_comb;
  wire [31:0] p7_add_63215_comb;
  wire [31:0] p7_add_63236_comb;
  wire [31:0] p7_add_63212_comb;
  wire [31:0] p7_add_63216_comb;
  wire [31:0] p7_add_63238_comb;
  assign p7_and_63217_comb = p6_add_63162 & p6_add_63084;
  assign p7_add_63210_comb = (p6_add_63134 & p6_add_63058 ^ ~(p6_add_63134 | ~p6_add_62982)) + {p6_add_63134[5:0] ^ p6_add_63134[10:5] ^ p6_add_63134[24:19], p6_add_63134[31:27] ^ p6_add_63134[4:0] ^ p6_add_63134[18:14], p6_add_63134[26:13] ^ p6_add_63134[31:18] ^ p6_add_63134[13:0], p6_add_63134[12:6] ^ p6_add_63134[17:11] ^ p6_add_63134[31:25]};
  assign p7_bit_slice_63213_comb = p6_message[287:256];
  assign p7_add_63211_comb = p7_add_63210_comb + p6_add_63140;
  assign p7_add_63215_comb = p7_bit_slice_63213_comb + 32'hab1c_5ed5;
  assign p7_add_63236_comb = (p7_and_63217_comb ^ p6_add_63162 & p6_add_63010 ^ p6_and_63141) + p6_add_63133;
  assign p7_add_63212_comb = p7_add_63211_comb + p6_add_63010;
  assign p7_add_63216_comb = p6_add_62982 + p7_add_63215_comb;
  assign p7_add_63238_comb = p7_add_63236_comb + {p6_add_63162[1:0] ^ p6_add_63162[12:11] ^ p6_add_63162[21:20], p6_add_63162[31:21] ^ p6_add_63162[10:0] ^ p6_add_63162[19:9], p6_add_63162[20:12] ^ p6_add_63162[31:23] ^ p6_add_63162[8:0], p6_add_63162[11:2] ^ p6_add_63162[22:13] ^ p6_add_63162[31:22]};

  // Registers for pipe stage 7:
  reg [511:0] p7_message;
  reg [31:0] p7_bit_slice_62886;
  reg [31:0] p7_bit_slice_62984;
  reg [31:0] p7_add_63058;
  reg [31:0] p7_bit_slice_63059;
  reg [31:0] p7_add_63134;
  reg [31:0] p7_add_63211;
  reg [31:0] p7_add_63212;
  reg [31:0] p7_bit_slice_63213;
  reg [31:0] p7_add_63216;
  reg [31:0] p7_add_63084;
  reg [31:0] p7_add_63162;
  reg [31:0] p7_and_63217;
  reg [31:0] p7_add_63238;
  always_ff @ (posedge clk) begin
    p7_message <= p6_message;
    p7_bit_slice_62886 <= p6_bit_slice_62886;
    p7_bit_slice_62984 <= p6_bit_slice_62984;
    p7_add_63058 <= p6_add_63058;
    p7_bit_slice_63059 <= p6_bit_slice_63059;
    p7_add_63134 <= p6_add_63134;
    p7_add_63211 <= p7_add_63211_comb;
    p7_add_63212 <= p7_add_63212_comb;
    p7_bit_slice_63213 <= p7_bit_slice_63213_comb;
    p7_add_63216 <= p7_add_63216_comb;
    p7_add_63084 <= p6_add_63084;
    p7_add_63162 <= p6_add_63162;
    p7_and_63217 <= p7_and_63217_comb;
    p7_add_63238 <= p7_add_63238_comb;
  end

  // ===== Pipe stage 8:
  wire [31:0] p8_and_63297_comb;
  wire [31:0] p8_add_63288_comb;
  wire [28:0] p8_add_63293_comb;
  wire [31:0] p8_add_63289_comb;
  wire [31:0] p8_add_63316_comb;
  wire [31:0] p8_add_63290_comb;
  wire [31:0] p8_add_63296_comb;
  wire [31:0] p8_add_63318_comb;
  assign p8_and_63297_comb = p7_add_63238 & p7_add_63162;
  assign p8_add_63288_comb = {p7_add_63212[5:0] ^ p7_add_63212[10:5] ^ p7_add_63212[24:19], p7_add_63212[31:27] ^ p7_add_63212[4:0] ^ p7_add_63212[18:14], p7_add_63212[26:13] ^ p7_add_63212[31:18] ^ p7_add_63212[13:0], p7_add_63212[12:6] ^ p7_add_63212[17:11] ^ p7_add_63212[31:25]} + (p7_add_63212 & p7_add_63134 ^ ~(p7_add_63212 | ~p7_add_63058));
  assign p8_add_63293_comb = p7_message[255:227] + 29'h1b00_f553;
  assign p8_add_63289_comb = p8_add_63288_comb + p7_add_63216;
  assign p8_add_63316_comb = (p8_and_63297_comb ^ p7_add_63238 & p7_add_63084 ^ p7_and_63217) + p7_add_63211;
  assign p8_add_63290_comb = p8_add_63289_comb + p7_add_63084;
  assign p8_add_63296_comb = {p8_add_63293_comb, p7_message[226:224]} + p7_add_63058;
  assign p8_add_63318_comb = p8_add_63316_comb + {p7_add_63238[1:0] ^ p7_add_63238[12:11] ^ p7_add_63238[21:20], p7_add_63238[31:21] ^ p7_add_63238[10:0] ^ p7_add_63238[19:9], p7_add_63238[20:12] ^ p7_add_63238[31:23] ^ p7_add_63238[8:0], p7_add_63238[11:2] ^ p7_add_63238[22:13] ^ p7_add_63238[31:22]};

  // Registers for pipe stage 8:
  reg [511:0] p8_message;
  reg [31:0] p8_bit_slice_62886;
  reg [31:0] p8_bit_slice_62984;
  reg [31:0] p8_bit_slice_63059;
  reg [31:0] p8_add_63134;
  reg [31:0] p8_add_63212;
  reg [31:0] p8_bit_slice_63213;
  reg [31:0] p8_add_63289;
  reg [31:0] p8_add_63290;
  reg [31:0] p8_add_63296;
  reg [31:0] p8_add_63162;
  reg [31:0] p8_add_63238;
  reg [31:0] p8_and_63297;
  reg [31:0] p8_add_63318;
  always_ff @ (posedge clk) begin
    p8_message <= p7_message;
    p8_bit_slice_62886 <= p7_bit_slice_62886;
    p8_bit_slice_62984 <= p7_bit_slice_62984;
    p8_bit_slice_63059 <= p7_bit_slice_63059;
    p8_add_63134 <= p7_add_63134;
    p8_add_63212 <= p7_add_63212;
    p8_bit_slice_63213 <= p7_bit_slice_63213;
    p8_add_63289 <= p8_add_63289_comb;
    p8_add_63290 <= p8_add_63290_comb;
    p8_add_63296 <= p8_add_63296_comb;
    p8_add_63162 <= p7_add_63162;
    p8_add_63238 <= p7_add_63238;
    p8_and_63297 <= p8_and_63297_comb;
    p8_add_63318 <= p8_add_63318_comb;
  end

  // ===== Pipe stage 9:
  wire [31:0] p9_bit_slice_63371_comb;
  wire [31:0] p9_add_63430_comb;
  wire [31:0] p9_add_63431_comb;
  wire [31:0] p9_add_63432_comb;
  wire [31:0] p9_and_63375_comb;
  wire [31:0] p9_add_63368_comb;
  wire [31:0] p9_add_63369_comb;
  wire [31:0] p9_add_63373_comb;
  wire [31:0] p9_add_63394_comb;
  wire [31:0] p9_add_63370_comb;
  wire [31:0] p9_add_63374_comb;
  wire [31:0] p9_add_63396_comb;
  wire [31:0] p9_add_63449_comb;
  assign p9_bit_slice_63371_comb = p8_message[223:192];
  assign p9_add_63430_comb = p9_bit_slice_63371_comb + {p8_message[454:452] ^ p8_message[465:463], p8_message[451:448] ^ p8_message[462:459] ^ p8_message[479:476], p8_message[479:469] ^ p8_message[458:448] ^ p8_message[475:465], p8_message[468:455] ^ p8_message[479:466] ^ p8_message[464:451]};
  assign p9_add_63431_comb = {p8_message[48:39] ^ p8_message[50:41], p8_message[38:32] ^ p8_message[40:34] ^ p8_message[63:57], p8_message[63:62] ^ p8_message[33:32] ^ p8_message[56:55], p8_message[61:49] ^ p8_message[63:51] ^ p8_message[54:42]} + p8_message[511:480];
  assign p9_add_63432_comb = p9_add_63430_comb + p9_add_63431_comb;
  assign p9_and_63375_comb = p8_add_63318 & p8_add_63238;
  assign p9_add_63368_comb = (p8_add_63290 & p8_add_63212 ^ ~(p8_add_63290 | ~p8_add_63134)) + {p8_add_63290[5:0] ^ p8_add_63290[10:5] ^ p8_add_63290[24:19], p8_add_63290[31:27] ^ p8_add_63290[4:0] ^ p8_add_63290[18:14], p8_add_63290[26:13] ^ p8_add_63290[31:18] ^ p8_add_63290[13:0], p8_add_63290[12:6] ^ p8_add_63290[17:11] ^ p8_add_63290[31:25]};
  assign p9_add_63369_comb = p9_add_63368_comb + p8_add_63296;
  assign p9_add_63373_comb = p9_bit_slice_63371_comb + 32'h1283_5b01;
  assign p9_add_63394_comb = (p9_and_63375_comb ^ p8_add_63318 & p8_add_63162 ^ p8_and_63297) + p8_add_63289;
  assign p9_add_63370_comb = p9_add_63369_comb + p8_add_63162;
  assign p9_add_63374_comb = p8_add_63134 + p9_add_63373_comb;
  assign p9_add_63396_comb = p9_add_63394_comb + {p8_add_63318[1:0] ^ p8_add_63318[12:11] ^ p8_add_63318[21:20], p8_add_63318[31:21] ^ p8_add_63318[10:0] ^ p8_add_63318[19:9], p8_add_63318[20:12] ^ p8_add_63318[31:23] ^ p8_add_63318[8:0], p8_add_63318[11:2] ^ p8_add_63318[22:13] ^ p8_add_63318[31:22]};
  assign p9_add_63449_comb = {p9_add_63432_comb[16:7] ^ p9_add_63432_comb[18:9], p9_add_63432_comb[6:0] ^ p9_add_63432_comb[8:2] ^ p9_add_63432_comb[31:25], p9_add_63432_comb[31:30] ^ p9_add_63432_comb[1:0] ^ p9_add_63432_comb[24:23], p9_add_63432_comb[29:17] ^ p9_add_63432_comb[31:19] ^ p9_add_63432_comb[22:10]} + p8_bit_slice_62886;

  // Registers for pipe stage 9:
  reg [511:0] p9_message;
  reg [31:0] p9_bit_slice_62984;
  reg [31:0] p9_bit_slice_63059;
  reg [31:0] p9_add_63212;
  reg [31:0] p9_bit_slice_63213;
  reg [31:0] p9_add_63290;
  reg [31:0] p9_add_63369;
  reg [31:0] p9_add_63370;
  reg [31:0] p9_bit_slice_63371;
  reg [31:0] p9_add_63374;
  reg [31:0] p9_add_63238;
  reg [31:0] p9_add_63318;
  reg [31:0] p9_and_63375;
  reg [31:0] p9_add_63396;
  reg [31:0] p9_add_63432;
  reg [31:0] p9_add_63449;
  always_ff @ (posedge clk) begin
    p9_message <= p8_message;
    p9_bit_slice_62984 <= p8_bit_slice_62984;
    p9_bit_slice_63059 <= p8_bit_slice_63059;
    p9_add_63212 <= p8_add_63212;
    p9_bit_slice_63213 <= p8_bit_slice_63213;
    p9_add_63290 <= p8_add_63290;
    p9_add_63369 <= p9_add_63369_comb;
    p9_add_63370 <= p9_add_63370_comb;
    p9_bit_slice_63371 <= p9_bit_slice_63371_comb;
    p9_add_63374 <= p9_add_63374_comb;
    p9_add_63238 <= p8_add_63238;
    p9_add_63318 <= p8_add_63318;
    p9_and_63375 <= p9_and_63375_comb;
    p9_add_63396 <= p9_add_63396_comb;
    p9_add_63432 <= p9_add_63432_comb;
    p9_add_63449 <= p9_add_63449_comb;
  end

  // ===== Pipe stage 10:
  wire [31:0] p10_bit_slice_63512_comb;
  wire [31:0] p10_add_63588_comb;
  wire [1:0] p10_bit_slice_63535_comb;
  wire [31:0] p10_add_63589_comb;
  wire [31:0] p10_and_63513_comb;
  wire [31:0] p10_add_63503_comb;
  wire [30:0] p10_add_63508_comb;
  wire [31:0] p10_bit_slice_63565_comb;
  wire [31:0] p10_add_63504_comb;
  wire [31:0] p10_add_63532_comb;
  wire [31:0] p10_add_63569_comb;
  wire [31:0] p10_add_63570_comb;
  wire [31:0] p10_bit_slice_63620_comb;
  wire [31:0] p10_add_63505_comb;
  wire [31:0] p10_add_63511_comb;
  wire [31:0] p10_add_63534_comb;
  wire [31:0] p10_add_63571_comb;
  wire [31:0] p10_add_63623_comb;
  wire [31:0] p10_add_63624_comb;
  assign p10_bit_slice_63512_comb = p9_message[159:128];
  assign p10_add_63588_comb = p10_bit_slice_63512_comb + {p9_message[390:388] ^ p9_message[401:399], p9_message[387:384] ^ p9_message[398:395] ^ p9_message[415:412], p9_message[415:405] ^ p9_message[394:384] ^ p9_message[411:401], p9_message[404:391] ^ p9_message[415:402] ^ p9_message[400:387]};
  assign p10_bit_slice_63535_comb = p9_message[1:0];
  assign p10_add_63589_comb = p10_add_63588_comb + p9_add_63449;
  assign p10_and_63513_comb = p9_add_63396 & p9_add_63318;
  assign p10_add_63503_comb = {p9_add_63370[5:0] ^ p9_add_63370[10:5] ^ p9_add_63370[24:19], p9_add_63370[31:27] ^ p9_add_63370[4:0] ^ p9_add_63370[18:14], p9_add_63370[26:13] ^ p9_add_63370[31:18] ^ p9_add_63370[13:0], p9_add_63370[12:6] ^ p9_add_63370[17:11] ^ p9_add_63370[31:25]} + (p9_add_63370 & p9_add_63290 ^ ~(p9_add_63370 | ~p9_add_63212));
  assign p10_add_63508_comb = p9_message[191:161] + 31'h1218_c2df;
  assign p10_bit_slice_63565_comb = p9_message[191:160];
  assign p10_add_63504_comb = p10_add_63503_comb + p9_add_63374;
  assign p10_add_63532_comb = (p10_and_63513_comb ^ p9_add_63396 & p9_add_63238 ^ p9_and_63375) + p9_add_63369;
  assign p10_add_63569_comb = p10_bit_slice_63565_comb + {p9_message[422:420] ^ p9_message[433:431], p9_message[419:416] ^ p9_message[430:427] ^ p9_message[447:444], p9_message[447:437] ^ p9_message[426:416] ^ p9_message[443:433], p9_message[436:423] ^ p9_message[447:434] ^ p9_message[432:419]};
  assign p10_add_63570_comb = {p9_message[16:7] ^ p9_message[18:9], p9_message[6:0] ^ p9_message[8:2] ^ p9_message[31:25], p9_message[31:30] ^ p10_bit_slice_63535_comb ^ p9_message[24:23], p9_message[29:17] ^ p9_message[31:19] ^ p9_message[22:10]} + p9_message[479:448];
  assign p10_bit_slice_63620_comb = p9_message[95:64];
  assign p10_add_63505_comb = p10_add_63504_comb + p9_add_63238;
  assign p10_add_63511_comb = {p10_add_63508_comb, p9_message[160]} + p9_add_63212;
  assign p10_add_63534_comb = p10_add_63532_comb + {p9_add_63396[1:0] ^ p9_add_63396[12:11] ^ p9_add_63396[21:20], p9_add_63396[31:21] ^ p9_add_63396[10:0] ^ p9_add_63396[19:9], p9_add_63396[20:12] ^ p9_add_63396[31:23] ^ p9_add_63396[8:0], p9_add_63396[11:2] ^ p9_add_63396[22:13] ^ p9_add_63396[31:22]};
  assign p10_add_63571_comb = p10_add_63569_comb + p10_add_63570_comb;
  assign p10_add_63623_comb = p10_bit_slice_63620_comb + {p9_message[326:324] ^ p9_message[337:335], p9_message[323:320] ^ p9_message[334:331] ^ p9_message[351:348], p9_message[351:341] ^ p9_message[330:320] ^ p9_message[347:337], p9_message[340:327] ^ p9_message[351:338] ^ p9_message[336:323]};
  assign p10_add_63624_comb = {p10_add_63589_comb[16:7] ^ p10_add_63589_comb[18:9], p10_add_63589_comb[6:0] ^ p10_add_63589_comb[8:2] ^ p10_add_63589_comb[31:25], p10_add_63589_comb[31:30] ^ p10_add_63589_comb[1:0] ^ p10_add_63589_comb[24:23], p10_add_63589_comb[29:17] ^ p10_add_63589_comb[31:19] ^ p10_add_63589_comb[22:10]} + p9_bit_slice_62984;

  // Registers for pipe stage 10:
  reg [511:0] p10_message;
  reg [31:0] p10_bit_slice_63059;
  reg [31:0] p10_bit_slice_63213;
  reg [31:0] p10_add_63290;
  reg [31:0] p10_add_63370;
  reg [31:0] p10_bit_slice_63371;
  reg [31:0] p10_add_63504;
  reg [31:0] p10_add_63505;
  reg [31:0] p10_add_63511;
  reg [31:0] p10_add_63318;
  reg [31:0] p10_bit_slice_63512;
  reg [31:0] p10_add_63396;
  reg [31:0] p10_and_63513;
  reg [31:0] p10_add_63534;
  reg [1:0] p10_bit_slice_63535;
  reg [31:0] p10_add_63432;
  reg [31:0] p10_bit_slice_63565;
  reg [31:0] p10_add_63571;
  reg [31:0] p10_add_63589;
  reg [31:0] p10_bit_slice_63620;
  reg [31:0] p10_add_63623;
  reg [31:0] p10_add_63624;
  always_ff @ (posedge clk) begin
    p10_message <= p9_message;
    p10_bit_slice_63059 <= p9_bit_slice_63059;
    p10_bit_slice_63213 <= p9_bit_slice_63213;
    p10_add_63290 <= p9_add_63290;
    p10_add_63370 <= p9_add_63370;
    p10_bit_slice_63371 <= p9_bit_slice_63371;
    p10_add_63504 <= p10_add_63504_comb;
    p10_add_63505 <= p10_add_63505_comb;
    p10_add_63511 <= p10_add_63511_comb;
    p10_add_63318 <= p9_add_63318;
    p10_bit_slice_63512 <= p10_bit_slice_63512_comb;
    p10_add_63396 <= p9_add_63396;
    p10_and_63513 <= p10_and_63513_comb;
    p10_add_63534 <= p10_add_63534_comb;
    p10_bit_slice_63535 <= p10_bit_slice_63535_comb;
    p10_add_63432 <= p9_add_63432;
    p10_bit_slice_63565 <= p10_bit_slice_63565_comb;
    p10_add_63571 <= p10_add_63571_comb;
    p10_add_63589 <= p10_add_63589_comb;
    p10_bit_slice_63620 <= p10_bit_slice_63620_comb;
    p10_add_63623 <= p10_add_63623_comb;
    p10_add_63624 <= p10_add_63624_comb;
  end

  // ===== Pipe stage 11:
  wire [31:0] p11_bit_slice_63767_comb;
  wire [31:0] p11_add_63771_comb;
  wire [31:0] p11_add_63772_comb;
  wire [31:0] p11_add_63775_comb;
  wire [31:0] p11_add_63773_comb;
  wire [31:0] p11_add_63690_comb;
  wire [31:0] p11_and_63708_comb;
  wire [1:0] p11_bit_slice_63774_comb;
  wire [31:0] p11_add_63691_comb;
  wire [29:0] p11_add_63700_comb;
  wire [30:0] p11_add_63706_comb;
  wire [31:0] p11_bit_slice_63839_comb;
  wire [31:0] p11_add_63692_comb;
  wire [31:0] p11_add_63696_comb;
  wire [31:0] p11_add_63729_comb;
  wire [29:0] p11_add_63735_comb;
  wire [31:0] p11_bit_slice_63732_comb;
  wire [31:0] p11_add_63843_comb;
  wire [31:0] p11_add_63844_comb;
  wire [31:0] p11_nor_63694_comb;
  wire [31:0] p11_add_63697_comb;
  wire [31:0] p11_add_63703_comb;
  wire [31:0] p11_add_63728_comb;
  wire [31:0] p11_add_63731_comb;
  wire [31:0] p11_concat_63736_comb;
  wire [31:0] p11_add_63807_comb;
  wire [31:0] p11_add_63808_comb;
  wire [31:0] p11_add_63845_comb;
  wire [31:0] p11_add_63862_comb;
  wire [31:0] p11_bit_slice_63879_comb;
  wire [31:0] p11_add_63880_comb;
  wire [31:0] p11_add_63897_comb;
  wire [31:0] p11_add_63914_comb;
  wire [31:0] p11_add_63931_comb;
  wire [31:0] p11_concat_63947_comb;
  wire [31:0] p11_concat_63963_comb;
  wire [31:0] p11_concat_63979_comb;
  assign p11_bit_slice_63767_comb = p10_message[127:96];
  assign p11_add_63771_comb = p11_bit_slice_63767_comb + {p10_message[358:356] ^ p10_message[369:367], p10_message[355:352] ^ p10_message[366:363] ^ p10_message[383:380], p10_message[383:373] ^ p10_message[362:352] ^ p10_message[379:369], p10_message[372:359] ^ p10_message[383:370] ^ p10_message[368:355]};
  assign p11_add_63772_comb = {p10_add_63571[16:7] ^ p10_add_63571[18:9], p10_add_63571[6:0] ^ p10_add_63571[8:2] ^ p10_add_63571[31:25], p10_add_63571[31:30] ^ p10_add_63571[1:0] ^ p10_add_63571[24:23], p10_add_63571[29:17] ^ p10_add_63571[31:19] ^ p10_add_63571[22:10]} + p10_message[415:384];
  assign p11_add_63775_comb = p10_add_63623 + p10_add_63624;
  assign p11_add_63773_comb = p11_add_63771_comb + p11_add_63772_comb;
  assign p11_add_63690_comb = (p10_add_63505 & p10_add_63370 ^ ~(p10_add_63505 | ~p10_add_63290)) + {p10_add_63505[5:0] ^ p10_add_63505[10:5] ^ p10_add_63505[24:19], p10_add_63505[31:27] ^ p10_add_63505[4:0] ^ p10_add_63505[18:14], p10_add_63505[26:13] ^ p10_add_63505[31:18] ^ p10_add_63505[13:0], p10_add_63505[12:6] ^ p10_add_63505[17:11] ^ p10_add_63505[31:25]};
  assign p11_and_63708_comb = p10_add_63534 & p10_add_63396;
  assign p11_bit_slice_63774_comb = p11_add_63773_comb[1:0];
  assign p11_add_63691_comb = p11_add_63690_comb + p10_add_63511;
  assign p11_add_63700_comb = p10_message[127:98] + 30'h1caf_975d;
  assign p11_add_63706_comb = p10_message[95:65] + 31'h406f_58ff;
  assign p11_bit_slice_63839_comb = p10_message[31:0];
  assign p11_add_63692_comb = p11_add_63691_comb + p10_add_63318;
  assign p11_add_63696_comb = p10_bit_slice_63512 + 32'h550c_7dc3;
  assign p11_add_63729_comb = (p11_and_63708_comb ^ p10_add_63534 & p10_add_63318 ^ p10_and_63513) + p10_add_63504;
  assign p11_add_63735_comb = p10_message[31:2] + 30'h3066_fc5d;
  assign p11_bit_slice_63732_comb = p10_message[63:32];
  assign p11_add_63843_comb = p11_bit_slice_63839_comb + {p10_message[262:260] ^ p10_message[273:271], p10_message[259:256] ^ p10_message[270:267] ^ p10_message[287:284], p10_message[287:277] ^ p10_message[266:256] ^ p10_message[283:273], p10_message[276:263] ^ p10_message[287:274] ^ p10_message[272:259]};
  assign p11_add_63844_comb = {p11_add_63775_comb[16:7] ^ p11_add_63775_comb[18:9], p11_add_63775_comb[6:0] ^ p11_add_63775_comb[8:2] ^ p11_add_63775_comb[31:25], p11_add_63775_comb[31:30] ^ p11_add_63775_comb[1:0] ^ p11_add_63775_comb[24:23], p11_add_63775_comb[29:17] ^ p11_add_63775_comb[31:19] ^ p11_add_63775_comb[22:10]} + p10_message[319:288];
  assign p11_nor_63694_comb = ~(p11_add_63692_comb | ~p10_add_63370);
  assign p11_add_63697_comb = p10_add_63290 + p11_add_63696_comb;
  assign p11_add_63703_comb = {p11_add_63700_comb, p10_message[97:96]} + p10_add_63370;
  assign p11_add_63728_comb = {p11_add_63706_comb, p10_message[64]} + p10_add_63505;
  assign p11_add_63731_comb = p11_add_63729_comb + {p10_add_63534[1:0] ^ p10_add_63534[12:11] ^ p10_add_63534[21:20], p10_add_63534[31:21] ^ p10_add_63534[10:0] ^ p10_add_63534[19:9], p10_add_63534[20:12] ^ p10_add_63534[31:23] ^ p10_add_63534[8:0], p10_add_63534[11:2] ^ p10_add_63534[22:13] ^ p10_add_63534[31:22]};
  assign p11_concat_63736_comb = {p11_add_63735_comb, p10_bit_slice_63535};
  assign p11_add_63807_comb = p11_bit_slice_63732_comb + {p10_message[294:292] ^ p10_message[305:303], p10_message[291:288] ^ p10_message[302:299] ^ p10_message[319:316], p10_message[319:309] ^ p10_message[298:288] ^ p10_message[315:305], p10_message[308:295] ^ p10_message[319:306] ^ p10_message[304:291]};
  assign p11_add_63808_comb = {p11_add_63773_comb[16:7] ^ p11_add_63773_comb[18:9], p11_add_63773_comb[6:0] ^ p11_add_63773_comb[8:2] ^ p11_add_63773_comb[31:25], p11_add_63773_comb[31:30] ^ p11_bit_slice_63774_comb ^ p11_add_63773_comb[24:23], p11_add_63773_comb[29:17] ^ p11_add_63773_comb[31:19] ^ p11_add_63773_comb[22:10]} + p10_bit_slice_63059;
  assign p11_add_63845_comb = p11_add_63843_comb + p11_add_63844_comb;
  assign p11_add_63862_comb = p10_add_63432 + {p10_message[230:228] ^ p10_message[241:239], p10_message[227:224] ^ p10_message[238:235] ^ p10_message[255:252], p10_message[255:245] ^ p10_message[234:224] ^ p10_message[251:241], p10_message[244:231] ^ p10_message[255:242] ^ p10_message[240:227]};
  assign p11_bit_slice_63879_comb = p10_message[255:224];
  assign p11_add_63880_comb = p10_add_63571 + {p10_message[198:196] ^ p10_message[209:207], p10_message[195:192] ^ p10_message[206:203] ^ p10_message[223:220], p10_message[223:213] ^ p10_message[202:192] ^ p10_message[219:209], p10_message[212:199] ^ p10_message[223:210] ^ p10_message[208:195]};
  assign p11_add_63897_comb = p10_add_63589 + {p10_message[166:164] ^ p10_message[177:175], p10_message[163:160] ^ p10_message[174:171] ^ p10_message[191:188], p10_message[191:181] ^ p10_message[170:160] ^ p10_message[187:177], p10_message[180:167] ^ p10_message[191:178] ^ p10_message[176:163]};
  assign p11_add_63914_comb = p11_add_63773_comb + {p10_message[134:132] ^ p10_message[145:143], p10_message[131:128] ^ p10_message[142:139] ^ p10_message[159:156], p10_message[159:149] ^ p10_message[138:128] ^ p10_message[155:145], p10_message[148:135] ^ p10_message[159:146] ^ p10_message[144:131]};
  assign p11_add_63931_comb = p11_add_63775_comb + {p10_message[102:100] ^ p10_message[113:111], p10_message[99:96] ^ p10_message[110:107] ^ p10_message[127:124], p10_message[127:117] ^ p10_message[106:96] ^ p10_message[123:113], p10_message[116:103] ^ p10_message[127:114] ^ p10_message[112:99]};
  assign p11_concat_63947_comb = {p10_message[70:68] ^ p10_message[81:79], p10_message[67:64] ^ p10_message[78:75] ^ p10_message[95:92], p10_message[95:85] ^ p10_message[74:64] ^ p10_message[91:81], p10_message[84:71] ^ p10_message[95:82] ^ p10_message[80:67]};
  assign p11_concat_63963_comb = {p10_message[38:36] ^ p10_message[49:47], p10_message[35:32] ^ p10_message[46:43] ^ p10_message[63:60], p10_message[63:53] ^ p10_message[42:32] ^ p10_message[59:49], p10_message[52:39] ^ p10_message[63:50] ^ p10_message[48:35]};
  assign p11_concat_63979_comb = {p10_message[6:4] ^ p10_message[17:15], p10_message[3:0] ^ p10_message[14:11] ^ p10_message[31:28], p10_message[31:21] ^ p10_message[10:0] ^ p10_message[27:17], p10_message[20:7] ^ p10_message[31:18] ^ p10_message[16:3]};

  // Registers for pipe stage 11:
  reg [31:0] p11_bit_slice_63213;
  reg [31:0] p11_bit_slice_63371;
  reg [31:0] p11_add_63505;
  reg [31:0] p11_add_63691;
  reg [31:0] p11_add_63692;
  reg [31:0] p11_nor_63694;
  reg [31:0] p11_bit_slice_63512;
  reg [31:0] p11_add_63697;
  reg [31:0] p11_add_63396;
  reg [31:0] p11_add_63703;
  reg [31:0] p11_add_63534;
  reg [31:0] p11_and_63708;
  reg [31:0] p11_add_63728;
  reg [31:0] p11_add_63731;
  reg [31:0] p11_bit_slice_63732;
  reg [31:0] p11_concat_63736;
  reg [31:0] p11_add_63432;
  reg [31:0] p11_bit_slice_63565;
  reg [31:0] p11_add_63571;
  reg [31:0] p11_add_63589;
  reg [31:0] p11_bit_slice_63767;
  reg [31:0] p11_add_63773;
  reg [1:0] p11_bit_slice_63774;
  reg [31:0] p11_bit_slice_63620;
  reg [31:0] p11_add_63775;
  reg [31:0] p11_add_63807;
  reg [31:0] p11_add_63808;
  reg [31:0] p11_bit_slice_63839;
  reg [31:0] p11_add_63845;
  reg [31:0] p11_add_63862;
  reg [31:0] p11_bit_slice_63879;
  reg [31:0] p11_add_63880;
  reg [31:0] p11_add_63897;
  reg [31:0] p11_add_63914;
  reg [31:0] p11_add_63931;
  reg [31:0] p11_concat_63947;
  reg [31:0] p11_concat_63963;
  reg [31:0] p11_concat_63979;
  always_ff @ (posedge clk) begin
    p11_bit_slice_63213 <= p10_bit_slice_63213;
    p11_bit_slice_63371 <= p10_bit_slice_63371;
    p11_add_63505 <= p10_add_63505;
    p11_add_63691 <= p11_add_63691_comb;
    p11_add_63692 <= p11_add_63692_comb;
    p11_nor_63694 <= p11_nor_63694_comb;
    p11_bit_slice_63512 <= p10_bit_slice_63512;
    p11_add_63697 <= p11_add_63697_comb;
    p11_add_63396 <= p10_add_63396;
    p11_add_63703 <= p11_add_63703_comb;
    p11_add_63534 <= p10_add_63534;
    p11_and_63708 <= p11_and_63708_comb;
    p11_add_63728 <= p11_add_63728_comb;
    p11_add_63731 <= p11_add_63731_comb;
    p11_bit_slice_63732 <= p11_bit_slice_63732_comb;
    p11_concat_63736 <= p11_concat_63736_comb;
    p11_add_63432 <= p10_add_63432;
    p11_bit_slice_63565 <= p10_bit_slice_63565;
    p11_add_63571 <= p10_add_63571;
    p11_add_63589 <= p10_add_63589;
    p11_bit_slice_63767 <= p11_bit_slice_63767_comb;
    p11_add_63773 <= p11_add_63773_comb;
    p11_bit_slice_63774 <= p11_bit_slice_63774_comb;
    p11_bit_slice_63620 <= p10_bit_slice_63620;
    p11_add_63775 <= p11_add_63775_comb;
    p11_add_63807 <= p11_add_63807_comb;
    p11_add_63808 <= p11_add_63808_comb;
    p11_bit_slice_63839 <= p11_bit_slice_63839_comb;
    p11_add_63845 <= p11_add_63845_comb;
    p11_add_63862 <= p11_add_63862_comb;
    p11_bit_slice_63879 <= p11_bit_slice_63879_comb;
    p11_add_63880 <= p11_add_63880_comb;
    p11_add_63897 <= p11_add_63897_comb;
    p11_add_63914 <= p11_add_63914_comb;
    p11_add_63931 <= p11_add_63931_comb;
    p11_concat_63947 <= p11_concat_63947_comb;
    p11_concat_63963 <= p11_concat_63963_comb;
    p11_concat_63979 <= p11_concat_63979_comb;
  end

  // ===== Pipe stage 12:
  wire [1:0] p12_bit_slice_64103_comb;
  wire [31:0] p12_add_64102_comb;
  wire [31:0] p12_add_64137_comb;
  wire [31:0] p12_add_64138_comb;
  wire [31:0] p12_add_64075_comb;
  wire [31:0] p12_and_64080_comb;
  wire [31:0] p12_add_64076_comb;
  wire [31:0] p12_add_64077_comb;
  wire [31:0] p12_add_64099_comb;
  wire [31:0] p12_add_64120_comb;
  wire [31:0] p12_nor_64079_comb;
  wire [31:0] p12_add_64101_comb;
  wire [31:0] p12_add_64121_comb;
  wire [31:0] p12_add_64155_comb;
  wire [31:0] p12_add_64156_comb;
  wire [31:0] p12_add_64157_comb;
  assign p12_bit_slice_64103_comb = p11_add_63845[1:0];
  assign p12_add_64102_comb = p11_add_63807 + p11_add_63808;
  assign p12_add_64137_comb = {p11_add_63845[16:7] ^ p11_add_63845[18:9], p11_add_63845[6:0] ^ p11_add_63845[8:2] ^ p11_add_63845[31:25], p11_add_63845[31:30] ^ p12_bit_slice_64103_comb ^ p11_add_63845[24:23], p11_add_63845[29:17] ^ p11_add_63845[31:19] ^ p11_add_63845[22:10]} + p11_bit_slice_63879;
  assign p12_add_64138_comb = p11_add_63880 + p12_add_64137_comb;
  assign p12_add_64075_comb = {p11_add_63692[5:0] ^ p11_add_63692[10:5] ^ p11_add_63692[24:19], p11_add_63692[31:27] ^ p11_add_63692[4:0] ^ p11_add_63692[18:14], p11_add_63692[26:13] ^ p11_add_63692[31:18] ^ p11_add_63692[13:0], p11_add_63692[12:6] ^ p11_add_63692[17:11] ^ p11_add_63692[31:25]} + (p11_add_63692 & p11_add_63505 ^ p11_nor_63694);
  assign p12_and_64080_comb = p11_add_63731 & p11_add_63534;
  assign p12_add_64076_comb = p12_add_64075_comb + p11_add_63697;
  assign p12_add_64077_comb = p12_add_64076_comb + p11_add_63396;
  assign p12_add_64099_comb = (p12_and_64080_comb ^ p11_add_63731 & p11_add_63396 ^ p11_and_63708) + p11_add_63691;
  assign p12_add_64120_comb = {p12_add_64102_comb[16:7] ^ p12_add_64102_comb[18:9], p12_add_64102_comb[6:0] ^ p12_add_64102_comb[8:2] ^ p12_add_64102_comb[31:25], p12_add_64102_comb[31:30] ^ p12_add_64102_comb[1:0] ^ p12_add_64102_comb[24:23], p12_add_64102_comb[29:17] ^ p12_add_64102_comb[31:19] ^ p12_add_64102_comb[22:10]} + p11_bit_slice_63213;
  assign p12_nor_64079_comb = ~(p12_add_64077_comb | ~p11_add_63505);
  assign p12_add_64101_comb = p12_add_64099_comb + {p11_add_63731[1:0] ^ p11_add_63731[12:11] ^ p11_add_63731[21:20], p11_add_63731[31:21] ^ p11_add_63731[10:0] ^ p11_add_63731[19:9], p11_add_63731[20:12] ^ p11_add_63731[31:23] ^ p11_add_63731[8:0], p11_add_63731[11:2] ^ p11_add_63731[22:13] ^ p11_add_63731[31:22]};
  assign p12_add_64121_comb = p11_add_63862 + p12_add_64120_comb;
  assign p12_add_64155_comb = {p12_add_64138_comb[16:7] ^ p12_add_64138_comb[18:9], p12_add_64138_comb[6:0] ^ p12_add_64138_comb[8:2] ^ p12_add_64138_comb[31:25], p12_add_64138_comb[31:30] ^ p12_add_64138_comb[1:0] ^ p12_add_64138_comb[24:23], p12_add_64138_comb[29:17] ^ p12_add_64138_comb[31:19] ^ p12_add_64138_comb[22:10]} + p11_bit_slice_63565;
  assign p12_add_64156_comb = p12_add_64102_comb + p11_concat_63947;
  assign p12_add_64157_comb = p11_add_63845 + p11_concat_63963;

  // Registers for pipe stage 12:
  reg [31:0] p12_bit_slice_63371;
  reg [31:0] p12_add_63692;
  reg [31:0] p12_bit_slice_63512;
  reg [31:0] p12_add_64076;
  reg [31:0] p12_add_64077;
  reg [31:0] p12_nor_64079;
  reg [31:0] p12_add_63703;
  reg [31:0] p12_add_63534;
  reg [31:0] p12_add_63728;
  reg [31:0] p12_add_63731;
  reg [31:0] p12_bit_slice_63732;
  reg [31:0] p12_and_64080;
  reg [31:0] p12_add_64101;
  reg [31:0] p12_concat_63736;
  reg [31:0] p12_add_63432;
  reg [31:0] p12_add_63571;
  reg [31:0] p12_add_63589;
  reg [31:0] p12_bit_slice_63767;
  reg [31:0] p12_add_63773;
  reg [1:0] p12_bit_slice_63774;
  reg [31:0] p12_bit_slice_63620;
  reg [31:0] p12_add_63775;
  reg [31:0] p12_add_64102;
  reg [31:0] p12_bit_slice_63839;
  reg [31:0] p12_add_63845;
  reg [1:0] p12_bit_slice_64103;
  reg [31:0] p12_add_64121;
  reg [31:0] p12_add_64138;
  reg [31:0] p12_add_63897;
  reg [31:0] p12_add_63914;
  reg [31:0] p12_add_64155;
  reg [31:0] p12_add_63931;
  reg [31:0] p12_add_64156;
  reg [31:0] p12_add_64157;
  reg [31:0] p12_concat_63979;
  always_ff @ (posedge clk) begin
    p12_bit_slice_63371 <= p11_bit_slice_63371;
    p12_add_63692 <= p11_add_63692;
    p12_bit_slice_63512 <= p11_bit_slice_63512;
    p12_add_64076 <= p12_add_64076_comb;
    p12_add_64077 <= p12_add_64077_comb;
    p12_nor_64079 <= p12_nor_64079_comb;
    p12_add_63703 <= p11_add_63703;
    p12_add_63534 <= p11_add_63534;
    p12_add_63728 <= p11_add_63728;
    p12_add_63731 <= p11_add_63731;
    p12_bit_slice_63732 <= p11_bit_slice_63732;
    p12_and_64080 <= p12_and_64080_comb;
    p12_add_64101 <= p12_add_64101_comb;
    p12_concat_63736 <= p11_concat_63736;
    p12_add_63432 <= p11_add_63432;
    p12_add_63571 <= p11_add_63571;
    p12_add_63589 <= p11_add_63589;
    p12_bit_slice_63767 <= p11_bit_slice_63767;
    p12_add_63773 <= p11_add_63773;
    p12_bit_slice_63774 <= p11_bit_slice_63774;
    p12_bit_slice_63620 <= p11_bit_slice_63620;
    p12_add_63775 <= p11_add_63775;
    p12_add_64102 <= p12_add_64102_comb;
    p12_bit_slice_63839 <= p11_bit_slice_63839;
    p12_add_63845 <= p11_add_63845;
    p12_bit_slice_64103 <= p12_bit_slice_64103_comb;
    p12_add_64121 <= p12_add_64121_comb;
    p12_add_64138 <= p12_add_64138_comb;
    p12_add_63897 <= p11_add_63897;
    p12_add_63914 <= p11_add_63914;
    p12_add_64155 <= p12_add_64155_comb;
    p12_add_63931 <= p11_add_63931;
    p12_add_64156 <= p12_add_64156_comb;
    p12_add_64157 <= p12_add_64157_comb;
    p12_concat_63979 <= p11_concat_63979;
  end

  // ===== Pipe stage 13:
  wire [31:0] p13_add_64289_comb;
  wire [31:0] p13_add_64291_comb;
  wire [31:0] p13_add_64290_comb;
  wire [31:0] p13_and_64250_comb;
  wire [31:0] p13_add_64247_comb;
  wire [31:0] p13_add_64248_comb;
  wire [31:0] p13_add_64270_comb;
  wire [31:0] p13_add_64325_comb;
  wire [31:0] p13_add_64249_comb;
  wire [31:0] p13_add_64269_comb;
  wire [31:0] p13_add_64272_comb;
  wire [31:0] p13_add_64308_comb;
  wire [31:0] p13_add_64326_comb;
  wire [31:0] p13_add_64327_comb;
  assign p13_add_64289_comb = {p12_add_64121[16:7] ^ p12_add_64121[18:9], p12_add_64121[6:0] ^ p12_add_64121[8:2] ^ p12_add_64121[31:25], p12_add_64121[31:30] ^ p12_add_64121[1:0] ^ p12_add_64121[24:23], p12_add_64121[29:17] ^ p12_add_64121[31:19] ^ p12_add_64121[22:10]} + p12_bit_slice_63371;
  assign p13_add_64291_comb = p12_add_63914 + p12_add_64155;
  assign p13_add_64290_comb = p12_add_63897 + p13_add_64289_comb;
  assign p13_and_64250_comb = p12_add_64101 & p12_add_63731;
  assign p13_add_64247_comb = (p12_add_64077 & p12_add_63692 ^ p12_nor_64079) + {p12_add_64077[5:0] ^ p12_add_64077[10:5] ^ p12_add_64077[24:19], p12_add_64077[31:27] ^ p12_add_64077[4:0] ^ p12_add_64077[18:14], p12_add_64077[26:13] ^ p12_add_64077[31:18] ^ p12_add_64077[13:0], p12_add_64077[12:6] ^ p12_add_64077[17:11] ^ p12_add_64077[31:25]};
  assign p13_add_64248_comb = p13_add_64247_comb + p12_add_63703;
  assign p13_add_64270_comb = (p13_and_64250_comb ^ p12_add_64101 & p12_add_63534 ^ p12_and_64080) + p12_add_64076;
  assign p13_add_64325_comb = {p13_add_64291_comb[16:7] ^ p13_add_64291_comb[18:9], p13_add_64291_comb[6:0] ^ p13_add_64291_comb[8:2] ^ p13_add_64291_comb[31:25], p13_add_64291_comb[31:30] ^ p13_add_64291_comb[1:0] ^ p13_add_64291_comb[24:23], p13_add_64291_comb[29:17] ^ p13_add_64291_comb[31:19] ^ p13_add_64291_comb[22:10]} + p12_bit_slice_63767;
  assign p13_add_64249_comb = p13_add_64248_comb + p12_add_63534;
  assign p13_add_64269_comb = p12_concat_63736 + p12_add_64077;
  assign p13_add_64272_comb = p13_add_64270_comb + {p12_add_64101[1:0] ^ p12_add_64101[12:11] ^ p12_add_64101[21:20], p12_add_64101[31:21] ^ p12_add_64101[10:0] ^ p12_add_64101[19:9], p12_add_64101[20:12] ^ p12_add_64101[31:23] ^ p12_add_64101[8:0], p12_add_64101[11:2] ^ p12_add_64101[22:13] ^ p12_add_64101[31:22]};
  assign p13_add_64308_comb = {p13_add_64290_comb[16:7] ^ p13_add_64290_comb[18:9], p13_add_64290_comb[6:0] ^ p13_add_64290_comb[8:2] ^ p13_add_64290_comb[31:25], p13_add_64290_comb[31:30] ^ p13_add_64290_comb[1:0] ^ p13_add_64290_comb[24:23], p13_add_64290_comb[29:17] ^ p13_add_64290_comb[31:19] ^ p13_add_64290_comb[22:10]} + p12_bit_slice_63512;
  assign p13_add_64326_comb = p12_add_64156 + p13_add_64325_comb;
  assign p13_add_64327_comb = p12_add_64121 + p12_concat_63979;

  // Registers for pipe stage 13:
  reg [31:0] p13_add_63692;
  reg [31:0] p13_add_64077;
  reg [31:0] p13_add_64248;
  reg [31:0] p13_add_64249;
  reg [31:0] p13_add_63728;
  reg [31:0] p13_add_63731;
  reg [31:0] p13_bit_slice_63732;
  reg [31:0] p13_add_64101;
  reg [31:0] p13_and_64250;
  reg [31:0] p13_add_64269;
  reg [31:0] p13_add_64272;
  reg [31:0] p13_add_63432;
  reg [31:0] p13_add_63571;
  reg [31:0] p13_add_63589;
  reg [31:0] p13_add_63773;
  reg [1:0] p13_bit_slice_63774;
  reg [31:0] p13_bit_slice_63620;
  reg [31:0] p13_add_63775;
  reg [31:0] p13_add_64102;
  reg [31:0] p13_bit_slice_63839;
  reg [31:0] p13_add_63845;
  reg [1:0] p13_bit_slice_64103;
  reg [31:0] p13_add_64121;
  reg [31:0] p13_add_64138;
  reg [31:0] p13_add_64290;
  reg [31:0] p13_add_64291;
  reg [31:0] p13_add_63931;
  reg [31:0] p13_add_64308;
  reg [31:0] p13_add_64326;
  reg [31:0] p13_add_64157;
  reg [31:0] p13_add_64327;
  always_ff @ (posedge clk) begin
    p13_add_63692 <= p12_add_63692;
    p13_add_64077 <= p12_add_64077;
    p13_add_64248 <= p13_add_64248_comb;
    p13_add_64249 <= p13_add_64249_comb;
    p13_add_63728 <= p12_add_63728;
    p13_add_63731 <= p12_add_63731;
    p13_bit_slice_63732 <= p12_bit_slice_63732;
    p13_add_64101 <= p12_add_64101;
    p13_and_64250 <= p13_and_64250_comb;
    p13_add_64269 <= p13_add_64269_comb;
    p13_add_64272 <= p13_add_64272_comb;
    p13_add_63432 <= p12_add_63432;
    p13_add_63571 <= p12_add_63571;
    p13_add_63589 <= p12_add_63589;
    p13_add_63773 <= p12_add_63773;
    p13_bit_slice_63774 <= p12_bit_slice_63774;
    p13_bit_slice_63620 <= p12_bit_slice_63620;
    p13_add_63775 <= p12_add_63775;
    p13_add_64102 <= p12_add_64102;
    p13_bit_slice_63839 <= p12_bit_slice_63839;
    p13_add_63845 <= p12_add_63845;
    p13_bit_slice_64103 <= p12_bit_slice_64103;
    p13_add_64121 <= p12_add_64121;
    p13_add_64138 <= p12_add_64138;
    p13_add_64290 <= p13_add_64290_comb;
    p13_add_64291 <= p13_add_64291_comb;
    p13_add_63931 <= p12_add_63931;
    p13_add_64308 <= p13_add_64308_comb;
    p13_add_64326 <= p13_add_64326_comb;
    p13_add_64157 <= p12_add_64157;
    p13_add_64327 <= p13_add_64327_comb;
  end

  // ===== Pipe stage 14:
  wire [31:0] p14_add_64441_comb;
  wire [31:0] p14_add_64411_comb;
  wire [31:0] p14_and_64419_comb;
  wire [31:0] p14_add_64412_comb;
  wire [31:0] p14_add_64413_comb;
  wire [31:0] p14_add_64417_comb;
  wire [31:0] p14_add_64438_comb;
  wire [31:0] p14_add_64458_comb;
  wire [31:0] p14_add_64476_comb;
  wire [31:0] p14_nor_64415_comb;
  wire [31:0] p14_add_64418_comb;
  wire [31:0] p14_add_64440_comb;
  wire [31:0] p14_add_64459_comb;
  wire [31:0] p14_add_64477_comb;
  assign p14_add_64441_comb = p13_add_63931 + p13_add_64308;
  assign p14_add_64411_comb = (p13_add_64249 & p13_add_64077 ^ ~(p13_add_64249 | ~p13_add_63692)) + {p13_add_64249[5:0] ^ p13_add_64249[10:5] ^ p13_add_64249[24:19], p13_add_64249[31:27] ^ p13_add_64249[4:0] ^ p13_add_64249[18:14], p13_add_64249[26:13] ^ p13_add_64249[31:18] ^ p13_add_64249[13:0], p13_add_64249[12:6] ^ p13_add_64249[17:11] ^ p13_add_64249[31:25]};
  assign p14_and_64419_comb = p13_add_64272 & p13_add_64101;
  assign p14_add_64412_comb = p14_add_64411_comb + p13_add_63728;
  assign p14_add_64413_comb = p14_add_64412_comb + p13_add_63731;
  assign p14_add_64417_comb = p13_bit_slice_63732 + 32'h9bdc_06a7;
  assign p14_add_64438_comb = (p14_and_64419_comb ^ p13_add_64272 & p13_add_63731 ^ p13_and_64250) + p13_add_64248;
  assign p14_add_64458_comb = {p14_add_64441_comb[16:7] ^ p14_add_64441_comb[18:9], p14_add_64441_comb[6:0] ^ p14_add_64441_comb[8:2] ^ p14_add_64441_comb[31:25], p14_add_64441_comb[31:30] ^ p14_add_64441_comb[1:0] ^ p14_add_64441_comb[24:23], p14_add_64441_comb[29:17] ^ p14_add_64441_comb[31:19] ^ p14_add_64441_comb[22:10]} + p13_bit_slice_63620;
  assign p14_add_64476_comb = {p13_add_64326[16:7] ^ p13_add_64326[18:9], p13_add_64326[6:0] ^ p13_add_64326[8:2] ^ p13_add_64326[31:25], p13_add_64326[31:30] ^ p13_add_64326[1:0] ^ p13_add_64326[24:23], p13_add_64326[29:17] ^ p13_add_64326[31:19] ^ p13_add_64326[22:10]} + p13_bit_slice_63732;
  assign p14_nor_64415_comb = ~(p14_add_64413_comb | ~p13_add_64077);
  assign p14_add_64418_comb = p13_add_63692 + p14_add_64417_comb;
  assign p14_add_64440_comb = p14_add_64438_comb + {p13_add_64272[1:0] ^ p13_add_64272[12:11] ^ p13_add_64272[21:20], p13_add_64272[31:21] ^ p13_add_64272[10:0] ^ p13_add_64272[19:9], p13_add_64272[20:12] ^ p13_add_64272[31:23] ^ p13_add_64272[8:0], p13_add_64272[11:2] ^ p13_add_64272[22:13] ^ p13_add_64272[31:22]};
  assign p14_add_64459_comb = p13_add_64157 + p14_add_64458_comb;
  assign p14_add_64477_comb = p13_add_64327 + p14_add_64476_comb;

  // Registers for pipe stage 14:
  reg [31:0] p14_add_64249;
  reg [31:0] p14_add_64412;
  reg [31:0] p14_add_64413;
  reg [31:0] p14_nor_64415;
  reg [31:0] p14_add_64418;
  reg [31:0] p14_add_64101;
  reg [31:0] p14_add_64269;
  reg [31:0] p14_add_64272;
  reg [31:0] p14_add_63432;
  reg [31:0] p14_and_64419;
  reg [31:0] p14_add_64440;
  reg [31:0] p14_add_63571;
  reg [31:0] p14_add_63589;
  reg [31:0] p14_add_63773;
  reg [1:0] p14_bit_slice_63774;
  reg [31:0] p14_add_63775;
  reg [31:0] p14_add_64102;
  reg [31:0] p14_bit_slice_63839;
  reg [31:0] p14_add_63845;
  reg [1:0] p14_bit_slice_64103;
  reg [31:0] p14_add_64121;
  reg [31:0] p14_add_64138;
  reg [31:0] p14_add_64290;
  reg [31:0] p14_add_64291;
  reg [31:0] p14_add_64441;
  reg [31:0] p14_add_64326;
  reg [31:0] p14_add_64459;
  reg [31:0] p14_add_64477;
  always_ff @ (posedge clk) begin
    p14_add_64249 <= p13_add_64249;
    p14_add_64412 <= p14_add_64412_comb;
    p14_add_64413 <= p14_add_64413_comb;
    p14_nor_64415 <= p14_nor_64415_comb;
    p14_add_64418 <= p14_add_64418_comb;
    p14_add_64101 <= p13_add_64101;
    p14_add_64269 <= p13_add_64269;
    p14_add_64272 <= p13_add_64272;
    p14_add_63432 <= p13_add_63432;
    p14_and_64419 <= p14_and_64419_comb;
    p14_add_64440 <= p14_add_64440_comb;
    p14_add_63571 <= p13_add_63571;
    p14_add_63589 <= p13_add_63589;
    p14_add_63773 <= p13_add_63773;
    p14_bit_slice_63774 <= p13_bit_slice_63774;
    p14_add_63775 <= p13_add_63775;
    p14_add_64102 <= p13_add_64102;
    p14_bit_slice_63839 <= p13_bit_slice_63839;
    p14_add_63845 <= p13_add_63845;
    p14_bit_slice_64103 <= p13_bit_slice_64103;
    p14_add_64121 <= p13_add_64121;
    p14_add_64138 <= p13_add_64138;
    p14_add_64290 <= p13_add_64290;
    p14_add_64291 <= p13_add_64291;
    p14_add_64441 <= p14_add_64441_comb;
    p14_add_64326 <= p13_add_64326;
    p14_add_64459 <= p14_add_64459_comb;
    p14_add_64477 <= p14_add_64477_comb;
  end

  // ===== Pipe stage 15:
  wire [31:0] p15_and_64556_comb;
  wire [31:0] p15_add_64553_comb;
  wire [31:0] p15_add_64554_comb;
  wire [31:0] p15_add_64575_comb;
  wire [31:0] p15_add_64610_comb;
  wire [31:0] p15_add_64611_comb;
  wire [31:0] p15_add_64555_comb;
  wire [31:0] p15_add_64577_comb;
  wire [31:0] p15_add_64612_comb;
  assign p15_and_64556_comb = p14_add_64440 & p14_add_64272;
  assign p15_add_64553_comb = {p14_add_64413[5:0] ^ p14_add_64413[10:5] ^ p14_add_64413[24:19], p14_add_64413[31:27] ^ p14_add_64413[4:0] ^ p14_add_64413[18:14], p14_add_64413[26:13] ^ p14_add_64413[31:18] ^ p14_add_64413[13:0], p14_add_64413[12:6] ^ p14_add_64413[17:11] ^ p14_add_64413[31:25]} + (p14_add_64413 & p14_add_64249 ^ p14_nor_64415);
  assign p15_add_64554_comb = p15_add_64553_comb + p14_add_64418;
  assign p15_add_64575_comb = (p15_and_64556_comb ^ p14_add_64440 & p14_add_64101 ^ p14_and_64419) + p14_add_64412;
  assign p15_add_64610_comb = p14_add_64138 + {p14_add_63432[6:4] ^ p14_add_63432[17:15], p14_add_63432[3:0] ^ p14_add_63432[14:11] ^ p14_add_63432[31:28], p14_add_63432[31:21] ^ p14_add_63432[10:0] ^ p14_add_63432[27:17], p14_add_63432[20:7] ^ p14_add_63432[31:18] ^ p14_add_63432[16:3]};
  assign p15_add_64611_comb = {p14_add_64459[16:7] ^ p14_add_64459[18:9], p14_add_64459[6:0] ^ p14_add_64459[8:2] ^ p14_add_64459[31:25], p14_add_64459[31:30] ^ p14_add_64459[1:0] ^ p14_add_64459[24:23], p14_add_64459[29:17] ^ p14_add_64459[31:19] ^ p14_add_64459[22:10]} + p14_bit_slice_63839;
  assign p15_add_64555_comb = p15_add_64554_comb + p14_add_64101;
  assign p15_add_64577_comb = p15_add_64575_comb + {p14_add_64440[1:0] ^ p14_add_64440[12:11] ^ p14_add_64440[21:20], p14_add_64440[31:21] ^ p14_add_64440[10:0] ^ p14_add_64440[19:9], p14_add_64440[20:12] ^ p14_add_64440[31:23] ^ p14_add_64440[8:0], p14_add_64440[11:2] ^ p14_add_64440[22:13] ^ p14_add_64440[31:22]};
  assign p15_add_64612_comb = p15_add_64610_comb + p15_add_64611_comb;

  // Registers for pipe stage 15:
  reg [31:0] p15_add_64249;
  reg [31:0] p15_add_64413;
  reg [31:0] p15_add_64554;
  reg [31:0] p15_add_64555;
  reg [31:0] p15_add_64269;
  reg [31:0] p15_add_64272;
  reg [31:0] p15_add_63432;
  reg [31:0] p15_add_64440;
  reg [31:0] p15_add_63571;
  reg [31:0] p15_and_64556;
  reg [31:0] p15_add_64577;
  reg [31:0] p15_add_63589;
  reg [31:0] p15_add_63773;
  reg [1:0] p15_bit_slice_63774;
  reg [31:0] p15_add_63775;
  reg [31:0] p15_add_64102;
  reg [31:0] p15_add_63845;
  reg [1:0] p15_bit_slice_64103;
  reg [31:0] p15_add_64121;
  reg [31:0] p15_add_64138;
  reg [31:0] p15_add_64290;
  reg [31:0] p15_add_64291;
  reg [31:0] p15_add_64441;
  reg [31:0] p15_add_64326;
  reg [31:0] p15_add_64459;
  reg [31:0] p15_add_64477;
  reg [31:0] p15_add_64612;
  always_ff @ (posedge clk) begin
    p15_add_64249 <= p14_add_64249;
    p15_add_64413 <= p14_add_64413;
    p15_add_64554 <= p15_add_64554_comb;
    p15_add_64555 <= p15_add_64555_comb;
    p15_add_64269 <= p14_add_64269;
    p15_add_64272 <= p14_add_64272;
    p15_add_63432 <= p14_add_63432;
    p15_add_64440 <= p14_add_64440;
    p15_add_63571 <= p14_add_63571;
    p15_and_64556 <= p15_and_64556_comb;
    p15_add_64577 <= p15_add_64577_comb;
    p15_add_63589 <= p14_add_63589;
    p15_add_63773 <= p14_add_63773;
    p15_bit_slice_63774 <= p14_bit_slice_63774;
    p15_add_63775 <= p14_add_63775;
    p15_add_64102 <= p14_add_64102;
    p15_add_63845 <= p14_add_63845;
    p15_bit_slice_64103 <= p14_bit_slice_64103;
    p15_add_64121 <= p14_add_64121;
    p15_add_64138 <= p14_add_64138;
    p15_add_64290 <= p14_add_64290;
    p15_add_64291 <= p14_add_64291;
    p15_add_64441 <= p14_add_64441;
    p15_add_64326 <= p14_add_64326;
    p15_add_64459 <= p14_add_64459;
    p15_add_64477 <= p14_add_64477;
    p15_add_64612 <= p15_add_64612_comb;
  end

  // ===== Pipe stage 16:
  wire [31:0] p16_and_64694_comb;
  wire [31:0] p16_add_64688_comb;
  wire [31:0] p16_add_64689_comb;
  wire [31:0] p16_add_64692_comb;
  wire [31:0] p16_add_64713_comb;
  wire [31:0] p16_add_64748_comb;
  wire [31:0] p16_add_64749_comb;
  wire [31:0] p16_add_64690_comb;
  wire [31:0] p16_add_64693_comb;
  wire [31:0] p16_add_64715_comb;
  wire [31:0] p16_add_64750_comb;
  assign p16_and_64694_comb = p15_add_64577 & p15_add_64440;
  assign p16_add_64688_comb = (p15_add_64555 & p15_add_64413 ^ ~(p15_add_64555 | ~p15_add_64249)) + {p15_add_64555[5:0] ^ p15_add_64555[10:5] ^ p15_add_64555[24:19], p15_add_64555[31:27] ^ p15_add_64555[4:0] ^ p15_add_64555[18:14], p15_add_64555[26:13] ^ p15_add_64555[31:18] ^ p15_add_64555[13:0], p15_add_64555[12:6] ^ p15_add_64555[17:11] ^ p15_add_64555[31:25]};
  assign p16_add_64689_comb = p16_add_64688_comb + p15_add_64269;
  assign p16_add_64692_comb = p15_add_63432 + 32'he49b_69c1;
  assign p16_add_64713_comb = (p16_and_64694_comb ^ p15_add_64577 & p15_add_64272 ^ p15_and_64556) + p15_add_64554;
  assign p16_add_64748_comb = p15_add_64290 + {p15_add_63571[6:4] ^ p15_add_63571[17:15], p15_add_63571[3:0] ^ p15_add_63571[14:11] ^ p15_add_63571[31:28], p15_add_63571[31:21] ^ p15_add_63571[10:0] ^ p15_add_63571[27:17], p15_add_63571[20:7] ^ p15_add_63571[31:18] ^ p15_add_63571[16:3]};
  assign p16_add_64749_comb = {p15_add_64477[16:7] ^ p15_add_64477[18:9], p15_add_64477[6:0] ^ p15_add_64477[8:2] ^ p15_add_64477[31:25], p15_add_64477[31:30] ^ p15_add_64477[1:0] ^ p15_add_64477[24:23], p15_add_64477[29:17] ^ p15_add_64477[31:19] ^ p15_add_64477[22:10]} + p15_add_63432;
  assign p16_add_64690_comb = p16_add_64689_comb + p15_add_64272;
  assign p16_add_64693_comb = p15_add_64249 + p16_add_64692_comb;
  assign p16_add_64715_comb = p16_add_64713_comb + {p15_add_64577[1:0] ^ p15_add_64577[12:11] ^ p15_add_64577[21:20], p15_add_64577[31:21] ^ p15_add_64577[10:0] ^ p15_add_64577[19:9], p15_add_64577[20:12] ^ p15_add_64577[31:23] ^ p15_add_64577[8:0], p15_add_64577[11:2] ^ p15_add_64577[22:13] ^ p15_add_64577[31:22]};
  assign p16_add_64750_comb = p16_add_64748_comb + p16_add_64749_comb;

  // Registers for pipe stage 16:
  reg [31:0] p16_add_64413;
  reg [31:0] p16_add_64555;
  reg [31:0] p16_add_64689;
  reg [31:0] p16_add_64690;
  reg [31:0] p16_add_64693;
  reg [31:0] p16_add_64440;
  reg [31:0] p16_add_63571;
  reg [31:0] p16_add_64577;
  reg [31:0] p16_add_63589;
  reg [31:0] p16_and_64694;
  reg [31:0] p16_add_64715;
  reg [31:0] p16_add_63773;
  reg [1:0] p16_bit_slice_63774;
  reg [31:0] p16_add_63775;
  reg [31:0] p16_add_64102;
  reg [31:0] p16_add_63845;
  reg [1:0] p16_bit_slice_64103;
  reg [31:0] p16_add_64121;
  reg [31:0] p16_add_64138;
  reg [31:0] p16_add_64290;
  reg [31:0] p16_add_64291;
  reg [31:0] p16_add_64441;
  reg [31:0] p16_add_64326;
  reg [31:0] p16_add_64459;
  reg [31:0] p16_add_64477;
  reg [31:0] p16_add_64612;
  reg [31:0] p16_add_64750;
  always_ff @ (posedge clk) begin
    p16_add_64413 <= p15_add_64413;
    p16_add_64555 <= p15_add_64555;
    p16_add_64689 <= p16_add_64689_comb;
    p16_add_64690 <= p16_add_64690_comb;
    p16_add_64693 <= p16_add_64693_comb;
    p16_add_64440 <= p15_add_64440;
    p16_add_63571 <= p15_add_63571;
    p16_add_64577 <= p15_add_64577;
    p16_add_63589 <= p15_add_63589;
    p16_and_64694 <= p16_and_64694_comb;
    p16_add_64715 <= p16_add_64715_comb;
    p16_add_63773 <= p15_add_63773;
    p16_bit_slice_63774 <= p15_bit_slice_63774;
    p16_add_63775 <= p15_add_63775;
    p16_add_64102 <= p15_add_64102;
    p16_add_63845 <= p15_add_63845;
    p16_bit_slice_64103 <= p15_bit_slice_64103;
    p16_add_64121 <= p15_add_64121;
    p16_add_64138 <= p15_add_64138;
    p16_add_64290 <= p15_add_64290;
    p16_add_64291 <= p15_add_64291;
    p16_add_64441 <= p15_add_64441;
    p16_add_64326 <= p15_add_64326;
    p16_add_64459 <= p15_add_64459;
    p16_add_64477 <= p15_add_64477;
    p16_add_64612 <= p15_add_64612;
    p16_add_64750 <= p16_add_64750_comb;
  end

  // ===== Pipe stage 17:
  wire [31:0] p17_and_64835_comb;
  wire [31:0] p17_add_64826_comb;
  wire [30:0] p17_add_64831_comb;
  wire [31:0] p17_add_64827_comb;
  wire [31:0] p17_add_64854_comb;
  wire [31:0] p17_add_64889_comb;
  wire [31:0] p17_add_64890_comb;
  wire [31:0] p17_add_64828_comb;
  wire [31:0] p17_add_64834_comb;
  wire [31:0] p17_add_64856_comb;
  wire [31:0] p17_add_64891_comb;
  assign p17_and_64835_comb = p16_add_64715 & p16_add_64577;
  assign p17_add_64826_comb = {p16_add_64690[5:0] ^ p16_add_64690[10:5] ^ p16_add_64690[24:19], p16_add_64690[31:27] ^ p16_add_64690[4:0] ^ p16_add_64690[18:14], p16_add_64690[26:13] ^ p16_add_64690[31:18] ^ p16_add_64690[13:0], p16_add_64690[12:6] ^ p16_add_64690[17:11] ^ p16_add_64690[31:25]} + (p16_add_64690 & p16_add_64555 ^ ~(p16_add_64690 | ~p16_add_64413));
  assign p17_add_64831_comb = p16_add_63571[31:1] + 31'h77df_23c3;
  assign p17_add_64827_comb = p17_add_64826_comb + p16_add_64693;
  assign p17_add_64854_comb = (p17_and_64835_comb ^ p16_add_64715 & p16_add_64440 ^ p16_and_64694) + p16_add_64689;
  assign p17_add_64889_comb = p16_add_64291 + {p16_add_63589[6:4] ^ p16_add_63589[17:15], p16_add_63589[3:0] ^ p16_add_63589[14:11] ^ p16_add_63589[31:28], p16_add_63589[31:21] ^ p16_add_63589[10:0] ^ p16_add_63589[27:17], p16_add_63589[20:7] ^ p16_add_63589[31:18] ^ p16_add_63589[16:3]};
  assign p17_add_64890_comb = {p16_add_64612[16:7] ^ p16_add_64612[18:9], p16_add_64612[6:0] ^ p16_add_64612[8:2] ^ p16_add_64612[31:25], p16_add_64612[31:30] ^ p16_add_64612[1:0] ^ p16_add_64612[24:23], p16_add_64612[29:17] ^ p16_add_64612[31:19] ^ p16_add_64612[22:10]} + p16_add_63571;
  assign p17_add_64828_comb = p17_add_64827_comb + p16_add_64440;
  assign p17_add_64834_comb = {p17_add_64831_comb, p16_add_63571[0]} + p16_add_64413;
  assign p17_add_64856_comb = p17_add_64854_comb + {p16_add_64715[1:0] ^ p16_add_64715[12:11] ^ p16_add_64715[21:20], p16_add_64715[31:21] ^ p16_add_64715[10:0] ^ p16_add_64715[19:9], p16_add_64715[20:12] ^ p16_add_64715[31:23] ^ p16_add_64715[8:0], p16_add_64715[11:2] ^ p16_add_64715[22:13] ^ p16_add_64715[31:22]};
  assign p17_add_64891_comb = p17_add_64889_comb + p17_add_64890_comb;

  // Registers for pipe stage 17:
  reg [31:0] p17_add_64555;
  reg [31:0] p17_add_64690;
  reg [31:0] p17_add_64827;
  reg [31:0] p17_add_64828;
  reg [31:0] p17_add_64834;
  reg [31:0] p17_add_64577;
  reg [31:0] p17_add_63589;
  reg [31:0] p17_add_64715;
  reg [31:0] p17_add_63773;
  reg [1:0] p17_bit_slice_63774;
  reg [31:0] p17_and_64835;
  reg [31:0] p17_add_64856;
  reg [31:0] p17_add_63775;
  reg [31:0] p17_add_64102;
  reg [31:0] p17_add_63845;
  reg [1:0] p17_bit_slice_64103;
  reg [31:0] p17_add_64121;
  reg [31:0] p17_add_64138;
  reg [31:0] p17_add_64290;
  reg [31:0] p17_add_64291;
  reg [31:0] p17_add_64441;
  reg [31:0] p17_add_64326;
  reg [31:0] p17_add_64459;
  reg [31:0] p17_add_64477;
  reg [31:0] p17_add_64612;
  reg [31:0] p17_add_64750;
  reg [31:0] p17_add_64891;
  always_ff @ (posedge clk) begin
    p17_add_64555 <= p16_add_64555;
    p17_add_64690 <= p16_add_64690;
    p17_add_64827 <= p17_add_64827_comb;
    p17_add_64828 <= p17_add_64828_comb;
    p17_add_64834 <= p17_add_64834_comb;
    p17_add_64577 <= p16_add_64577;
    p17_add_63589 <= p16_add_63589;
    p17_add_64715 <= p16_add_64715;
    p17_add_63773 <= p16_add_63773;
    p17_bit_slice_63774 <= p16_bit_slice_63774;
    p17_and_64835 <= p17_and_64835_comb;
    p17_add_64856 <= p17_add_64856_comb;
    p17_add_63775 <= p16_add_63775;
    p17_add_64102 <= p16_add_64102;
    p17_add_63845 <= p16_add_63845;
    p17_bit_slice_64103 <= p16_bit_slice_64103;
    p17_add_64121 <= p16_add_64121;
    p17_add_64138 <= p16_add_64138;
    p17_add_64290 <= p16_add_64290;
    p17_add_64291 <= p16_add_64291;
    p17_add_64441 <= p16_add_64441;
    p17_add_64326 <= p16_add_64326;
    p17_add_64459 <= p16_add_64459;
    p17_add_64477 <= p16_add_64477;
    p17_add_64612 <= p16_add_64612;
    p17_add_64750 <= p16_add_64750;
    p17_add_64891 <= p17_add_64891_comb;
  end

  // ===== Pipe stage 18:
  wire [31:0] p18_and_64976_comb;
  wire [31:0] p18_add_64967_comb;
  wire [30:0] p18_add_64972_comb;
  wire [31:0] p18_add_64968_comb;
  wire [31:0] p18_add_64995_comb;
  wire [31:0] p18_add_65030_comb;
  wire [31:0] p18_add_65031_comb;
  wire [31:0] p18_add_64969_comb;
  wire [31:0] p18_add_64975_comb;
  wire [31:0] p18_add_64997_comb;
  wire [31:0] p18_add_65032_comb;
  assign p18_and_64976_comb = p17_add_64856 & p17_add_64715;
  assign p18_add_64967_comb = (p17_add_64828 & p17_add_64690 ^ ~(p17_add_64828 | ~p17_add_64555)) + {p17_add_64828[5:0] ^ p17_add_64828[10:5] ^ p17_add_64828[24:19], p17_add_64828[31:27] ^ p17_add_64828[4:0] ^ p17_add_64828[18:14], p17_add_64828[26:13] ^ p17_add_64828[31:18] ^ p17_add_64828[13:0], p17_add_64828[12:6] ^ p17_add_64828[17:11] ^ p17_add_64828[31:25]};
  assign p18_add_64972_comb = p17_add_63589[31:1] + 31'h07e0_cee3;
  assign p18_add_64968_comb = p18_add_64967_comb + p17_add_64834;
  assign p18_add_64995_comb = (p18_and_64976_comb ^ p17_add_64856 & p17_add_64577 ^ p17_and_64835) + p17_add_64827;
  assign p18_add_65030_comb = p17_add_64441 + {p17_add_63773[6:4] ^ p17_add_63773[17:15], p17_add_63773[3:0] ^ p17_add_63773[14:11] ^ p17_add_63773[31:28], p17_add_63773[31:21] ^ p17_add_63773[10:0] ^ p17_add_63773[27:17], p17_add_63773[20:7] ^ p17_add_63773[31:18] ^ p17_add_63773[16:3]};
  assign p18_add_65031_comb = {p17_add_64750[16:7] ^ p17_add_64750[18:9], p17_add_64750[6:0] ^ p17_add_64750[8:2] ^ p17_add_64750[31:25], p17_add_64750[31:30] ^ p17_add_64750[1:0] ^ p17_add_64750[24:23], p17_add_64750[29:17] ^ p17_add_64750[31:19] ^ p17_add_64750[22:10]} + p17_add_63589;
  assign p18_add_64969_comb = p18_add_64968_comb + p17_add_64577;
  assign p18_add_64975_comb = {p18_add_64972_comb, p17_add_63589[0]} + p17_add_64555;
  assign p18_add_64997_comb = p18_add_64995_comb + {p17_add_64856[1:0] ^ p17_add_64856[12:11] ^ p17_add_64856[21:20], p17_add_64856[31:21] ^ p17_add_64856[10:0] ^ p17_add_64856[19:9], p17_add_64856[20:12] ^ p17_add_64856[31:23] ^ p17_add_64856[8:0], p17_add_64856[11:2] ^ p17_add_64856[22:13] ^ p17_add_64856[31:22]};
  assign p18_add_65032_comb = p18_add_65030_comb + p18_add_65031_comb;

  // Registers for pipe stage 18:
  reg [31:0] p18_add_64690;
  reg [31:0] p18_add_64828;
  reg [31:0] p18_add_64968;
  reg [31:0] p18_add_64969;
  reg [31:0] p18_add_64975;
  reg [31:0] p18_add_64715;
  reg [31:0] p18_add_63773;
  reg [1:0] p18_bit_slice_63774;
  reg [31:0] p18_add_64856;
  reg [31:0] p18_add_63775;
  reg [31:0] p18_and_64976;
  reg [31:0] p18_add_64997;
  reg [31:0] p18_add_64102;
  reg [31:0] p18_add_63845;
  reg [1:0] p18_bit_slice_64103;
  reg [31:0] p18_add_64121;
  reg [31:0] p18_add_64138;
  reg [31:0] p18_add_64290;
  reg [31:0] p18_add_64291;
  reg [31:0] p18_add_64441;
  reg [31:0] p18_add_64326;
  reg [31:0] p18_add_64459;
  reg [31:0] p18_add_64477;
  reg [31:0] p18_add_64612;
  reg [31:0] p18_add_64750;
  reg [31:0] p18_add_64891;
  reg [31:0] p18_add_65032;
  always_ff @ (posedge clk) begin
    p18_add_64690 <= p17_add_64690;
    p18_add_64828 <= p17_add_64828;
    p18_add_64968 <= p18_add_64968_comb;
    p18_add_64969 <= p18_add_64969_comb;
    p18_add_64975 <= p18_add_64975_comb;
    p18_add_64715 <= p17_add_64715;
    p18_add_63773 <= p17_add_63773;
    p18_bit_slice_63774 <= p17_bit_slice_63774;
    p18_add_64856 <= p17_add_64856;
    p18_add_63775 <= p17_add_63775;
    p18_and_64976 <= p18_and_64976_comb;
    p18_add_64997 <= p18_add_64997_comb;
    p18_add_64102 <= p17_add_64102;
    p18_add_63845 <= p17_add_63845;
    p18_bit_slice_64103 <= p17_bit_slice_64103;
    p18_add_64121 <= p17_add_64121;
    p18_add_64138 <= p17_add_64138;
    p18_add_64290 <= p17_add_64290;
    p18_add_64291 <= p17_add_64291;
    p18_add_64441 <= p17_add_64441;
    p18_add_64326 <= p17_add_64326;
    p18_add_64459 <= p17_add_64459;
    p18_add_64477 <= p17_add_64477;
    p18_add_64612 <= p17_add_64612;
    p18_add_64750 <= p17_add_64750;
    p18_add_64891 <= p17_add_64891;
    p18_add_65032 <= p18_add_65032_comb;
  end

  // ===== Pipe stage 19:
  wire [31:0] p19_and_65116_comb;
  wire [31:0] p19_add_65108_comb;
  wire [29:0] p19_add_65113_comb;
  wire [31:0] p19_add_65109_comb;
  wire [31:0] p19_add_65135_comb;
  wire [31:0] p19_add_65170_comb;
  wire [31:0] p19_add_65171_comb;
  wire [31:0] p19_add_65110_comb;
  wire [31:0] p19_add_65115_comb;
  wire [31:0] p19_add_65137_comb;
  wire [31:0] p19_add_65172_comb;
  assign p19_and_65116_comb = p18_add_64997 & p18_add_64856;
  assign p19_add_65108_comb = (p18_add_64969 & p18_add_64828 ^ ~(p18_add_64969 | ~p18_add_64690)) + {p18_add_64969[5:0] ^ p18_add_64969[10:5] ^ p18_add_64969[24:19], p18_add_64969[31:27] ^ p18_add_64969[4:0] ^ p18_add_64969[18:14], p18_add_64969[26:13] ^ p18_add_64969[31:18] ^ p18_add_64969[13:0], p18_add_64969[12:6] ^ p18_add_64969[17:11] ^ p18_add_64969[31:25]};
  assign p19_add_65113_comb = p18_add_63773[31:2] + 30'h0903_2873;
  assign p19_add_65109_comb = p19_add_65108_comb + p18_add_64975;
  assign p19_add_65135_comb = (p19_and_65116_comb ^ p18_add_64997 & p18_add_64715 ^ p18_and_64976) + p18_add_64968;
  assign p19_add_65170_comb = p18_add_64326 + {p18_add_63775[6:4] ^ p18_add_63775[17:15], p18_add_63775[3:0] ^ p18_add_63775[14:11] ^ p18_add_63775[31:28], p18_add_63775[31:21] ^ p18_add_63775[10:0] ^ p18_add_63775[27:17], p18_add_63775[20:7] ^ p18_add_63775[31:18] ^ p18_add_63775[16:3]};
  assign p19_add_65171_comb = {p18_add_64891[16:7] ^ p18_add_64891[18:9], p18_add_64891[6:0] ^ p18_add_64891[8:2] ^ p18_add_64891[31:25], p18_add_64891[31:30] ^ p18_add_64891[1:0] ^ p18_add_64891[24:23], p18_add_64891[29:17] ^ p18_add_64891[31:19] ^ p18_add_64891[22:10]} + p18_add_63773;
  assign p19_add_65110_comb = p19_add_65109_comb + p18_add_64715;
  assign p19_add_65115_comb = {p19_add_65113_comb, p18_bit_slice_63774} + p18_add_64690;
  assign p19_add_65137_comb = p19_add_65135_comb + {p18_add_64997[1:0] ^ p18_add_64997[12:11] ^ p18_add_64997[21:20], p18_add_64997[31:21] ^ p18_add_64997[10:0] ^ p18_add_64997[19:9], p18_add_64997[20:12] ^ p18_add_64997[31:23] ^ p18_add_64997[8:0], p18_add_64997[11:2] ^ p18_add_64997[22:13] ^ p18_add_64997[31:22]};
  assign p19_add_65172_comb = p19_add_65170_comb + p19_add_65171_comb;

  // Registers for pipe stage 19:
  reg [31:0] p19_add_64828;
  reg [31:0] p19_add_64969;
  reg [31:0] p19_add_65109;
  reg [31:0] p19_add_65110;
  reg [31:0] p19_add_65115;
  reg [31:0] p19_add_64856;
  reg [31:0] p19_add_63775;
  reg [31:0] p19_add_64997;
  reg [31:0] p19_add_64102;
  reg [31:0] p19_and_65116;
  reg [31:0] p19_add_65137;
  reg [31:0] p19_add_63845;
  reg [1:0] p19_bit_slice_64103;
  reg [31:0] p19_add_64121;
  reg [31:0] p19_add_64138;
  reg [31:0] p19_add_64290;
  reg [31:0] p19_add_64291;
  reg [31:0] p19_add_64441;
  reg [31:0] p19_add_64326;
  reg [31:0] p19_add_64459;
  reg [31:0] p19_add_64477;
  reg [31:0] p19_add_64612;
  reg [31:0] p19_add_64750;
  reg [31:0] p19_add_64891;
  reg [31:0] p19_add_65032;
  reg [31:0] p19_add_65172;
  always_ff @ (posedge clk) begin
    p19_add_64828 <= p18_add_64828;
    p19_add_64969 <= p18_add_64969;
    p19_add_65109 <= p19_add_65109_comb;
    p19_add_65110 <= p19_add_65110_comb;
    p19_add_65115 <= p19_add_65115_comb;
    p19_add_64856 <= p18_add_64856;
    p19_add_63775 <= p18_add_63775;
    p19_add_64997 <= p18_add_64997;
    p19_add_64102 <= p18_add_64102;
    p19_and_65116 <= p19_and_65116_comb;
    p19_add_65137 <= p19_add_65137_comb;
    p19_add_63845 <= p18_add_63845;
    p19_bit_slice_64103 <= p18_bit_slice_64103;
    p19_add_64121 <= p18_add_64121;
    p19_add_64138 <= p18_add_64138;
    p19_add_64290 <= p18_add_64290;
    p19_add_64291 <= p18_add_64291;
    p19_add_64441 <= p18_add_64441;
    p19_add_64326 <= p18_add_64326;
    p19_add_64459 <= p18_add_64459;
    p19_add_64477 <= p18_add_64477;
    p19_add_64612 <= p18_add_64612;
    p19_add_64750 <= p18_add_64750;
    p19_add_64891 <= p18_add_64891;
    p19_add_65032 <= p18_add_65032;
    p19_add_65172 <= p19_add_65172_comb;
  end

  // ===== Pipe stage 20:
  wire [31:0] p20_and_65252_comb;
  wire [31:0] p20_add_65246_comb;
  wire [31:0] p20_add_65247_comb;
  wire [31:0] p20_add_65250_comb;
  wire [31:0] p20_add_65271_comb;
  wire [31:0] p20_add_65248_comb;
  wire [31:0] p20_add_65251_comb;
  wire [31:0] p20_add_65273_comb;
  assign p20_and_65252_comb = p19_add_65137 & p19_add_64997;
  assign p20_add_65246_comb = (p19_add_65110 & p19_add_64969 ^ ~(p19_add_65110 | ~p19_add_64828)) + {p19_add_65110[5:0] ^ p19_add_65110[10:5] ^ p19_add_65110[24:19], p19_add_65110[31:27] ^ p19_add_65110[4:0] ^ p19_add_65110[18:14], p19_add_65110[26:13] ^ p19_add_65110[31:18] ^ p19_add_65110[13:0], p19_add_65110[12:6] ^ p19_add_65110[17:11] ^ p19_add_65110[31:25]};
  assign p20_add_65247_comb = p20_add_65246_comb + p19_add_65115;
  assign p20_add_65250_comb = p19_add_63775 + 32'h2de9_2c6f;
  assign p20_add_65271_comb = (p20_and_65252_comb ^ p19_add_65137 & p19_add_64856 ^ p19_and_65116) + p19_add_65109;
  assign p20_add_65248_comb = p20_add_65247_comb + p19_add_64856;
  assign p20_add_65251_comb = p19_add_64828 + p20_add_65250_comb;
  assign p20_add_65273_comb = p20_add_65271_comb + {p19_add_65137[1:0] ^ p19_add_65137[12:11] ^ p19_add_65137[21:20], p19_add_65137[31:21] ^ p19_add_65137[10:0] ^ p19_add_65137[19:9], p19_add_65137[20:12] ^ p19_add_65137[31:23] ^ p19_add_65137[8:0], p19_add_65137[11:2] ^ p19_add_65137[22:13] ^ p19_add_65137[31:22]};

  // Registers for pipe stage 20:
  reg [31:0] p20_add_64969;
  reg [31:0] p20_add_65110;
  reg [31:0] p20_add_65247;
  reg [31:0] p20_add_65248;
  reg [31:0] p20_add_63775;
  reg [31:0] p20_add_65251;
  reg [31:0] p20_add_64997;
  reg [31:0] p20_add_64102;
  reg [31:0] p20_add_65137;
  reg [31:0] p20_add_63845;
  reg [1:0] p20_bit_slice_64103;
  reg [31:0] p20_and_65252;
  reg [31:0] p20_add_65273;
  reg [31:0] p20_add_64121;
  reg [31:0] p20_add_64138;
  reg [31:0] p20_add_64290;
  reg [31:0] p20_add_64291;
  reg [31:0] p20_add_64441;
  reg [31:0] p20_add_64326;
  reg [31:0] p20_add_64459;
  reg [31:0] p20_add_64477;
  reg [31:0] p20_add_64612;
  reg [31:0] p20_add_64750;
  reg [31:0] p20_add_64891;
  reg [31:0] p20_add_65032;
  reg [31:0] p20_add_65172;
  always_ff @ (posedge clk) begin
    p20_add_64969 <= p19_add_64969;
    p20_add_65110 <= p19_add_65110;
    p20_add_65247 <= p20_add_65247_comb;
    p20_add_65248 <= p20_add_65248_comb;
    p20_add_63775 <= p19_add_63775;
    p20_add_65251 <= p20_add_65251_comb;
    p20_add_64997 <= p19_add_64997;
    p20_add_64102 <= p19_add_64102;
    p20_add_65137 <= p19_add_65137;
    p20_add_63845 <= p19_add_63845;
    p20_bit_slice_64103 <= p19_bit_slice_64103;
    p20_and_65252 <= p20_and_65252_comb;
    p20_add_65273 <= p20_add_65273_comb;
    p20_add_64121 <= p19_add_64121;
    p20_add_64138 <= p19_add_64138;
    p20_add_64290 <= p19_add_64290;
    p20_add_64291 <= p19_add_64291;
    p20_add_64441 <= p19_add_64441;
    p20_add_64326 <= p19_add_64326;
    p20_add_64459 <= p19_add_64459;
    p20_add_64477 <= p19_add_64477;
    p20_add_64612 <= p19_add_64612;
    p20_add_64750 <= p19_add_64750;
    p20_add_64891 <= p19_add_64891;
    p20_add_65032 <= p19_add_65032;
    p20_add_65172 <= p19_add_65172;
  end

  // ===== Pipe stage 21:
  wire [31:0] p21_and_65356_comb;
  wire [31:0] p21_add_65347_comb;
  wire [30:0] p21_add_65352_comb;
  wire [31:0] p21_add_65348_comb;
  wire [31:0] p21_add_65375_comb;
  wire [31:0] p21_add_65349_comb;
  wire [31:0] p21_add_65355_comb;
  wire [31:0] p21_add_65377_comb;
  assign p21_and_65356_comb = p20_add_65273 & p20_add_65137;
  assign p21_add_65347_comb = {p20_add_65248[5:0] ^ p20_add_65248[10:5] ^ p20_add_65248[24:19], p20_add_65248[31:27] ^ p20_add_65248[4:0] ^ p20_add_65248[18:14], p20_add_65248[26:13] ^ p20_add_65248[31:18] ^ p20_add_65248[13:0], p20_add_65248[12:6] ^ p20_add_65248[17:11] ^ p20_add_65248[31:25]} + (p20_add_65248 & p20_add_65110 ^ ~(p20_add_65248 | ~p20_add_64969));
  assign p21_add_65352_comb = p20_add_64102[31:1] + 31'h253a_4255;
  assign p21_add_65348_comb = p21_add_65347_comb + p20_add_65251;
  assign p21_add_65375_comb = (p21_and_65356_comb ^ p20_add_65273 & p20_add_64997 ^ p20_and_65252) + p20_add_65247;
  assign p21_add_65349_comb = p21_add_65348_comb + p20_add_64997;
  assign p21_add_65355_comb = {p21_add_65352_comb, p20_add_64102[0]} + p20_add_64969;
  assign p21_add_65377_comb = p21_add_65375_comb + {p20_add_65273[1:0] ^ p20_add_65273[12:11] ^ p20_add_65273[21:20], p20_add_65273[31:21] ^ p20_add_65273[10:0] ^ p20_add_65273[19:9], p20_add_65273[20:12] ^ p20_add_65273[31:23] ^ p20_add_65273[8:0], p20_add_65273[11:2] ^ p20_add_65273[22:13] ^ p20_add_65273[31:22]};

  // Registers for pipe stage 21:
  reg [31:0] p21_add_65110;
  reg [31:0] p21_add_65248;
  reg [31:0] p21_add_63775;
  reg [31:0] p21_add_65348;
  reg [31:0] p21_add_65349;
  reg [31:0] p21_add_64102;
  reg [31:0] p21_add_65355;
  reg [31:0] p21_add_65137;
  reg [31:0] p21_add_63845;
  reg [1:0] p21_bit_slice_64103;
  reg [31:0] p21_add_65273;
  reg [31:0] p21_add_64121;
  reg [31:0] p21_and_65356;
  reg [31:0] p21_add_65377;
  reg [31:0] p21_add_64138;
  reg [31:0] p21_add_64290;
  reg [31:0] p21_add_64291;
  reg [31:0] p21_add_64441;
  reg [31:0] p21_add_64326;
  reg [31:0] p21_add_64459;
  reg [31:0] p21_add_64477;
  reg [31:0] p21_add_64612;
  reg [31:0] p21_add_64750;
  reg [31:0] p21_add_64891;
  reg [31:0] p21_add_65032;
  reg [31:0] p21_add_65172;
  always_ff @ (posedge clk) begin
    p21_add_65110 <= p20_add_65110;
    p21_add_65248 <= p20_add_65248;
    p21_add_63775 <= p20_add_63775;
    p21_add_65348 <= p21_add_65348_comb;
    p21_add_65349 <= p21_add_65349_comb;
    p21_add_64102 <= p20_add_64102;
    p21_add_65355 <= p21_add_65355_comb;
    p21_add_65137 <= p20_add_65137;
    p21_add_63845 <= p20_add_63845;
    p21_bit_slice_64103 <= p20_bit_slice_64103;
    p21_add_65273 <= p20_add_65273;
    p21_add_64121 <= p20_add_64121;
    p21_and_65356 <= p21_and_65356_comb;
    p21_add_65377 <= p21_add_65377_comb;
    p21_add_64138 <= p20_add_64138;
    p21_add_64290 <= p20_add_64290;
    p21_add_64291 <= p20_add_64291;
    p21_add_64441 <= p20_add_64441;
    p21_add_64326 <= p20_add_64326;
    p21_add_64459 <= p20_add_64459;
    p21_add_64477 <= p20_add_64477;
    p21_add_64612 <= p20_add_64612;
    p21_add_64750 <= p20_add_64750;
    p21_add_64891 <= p20_add_64891;
    p21_add_65032 <= p20_add_65032;
    p21_add_65172 <= p20_add_65172;
  end

  // ===== Pipe stage 22:
  wire [31:0] p22_and_65459_comb;
  wire [31:0] p22_add_65451_comb;
  wire [29:0] p22_add_65456_comb;
  wire [31:0] p22_add_65452_comb;
  wire [31:0] p22_add_65478_comb;
  wire [31:0] p22_add_65453_comb;
  wire [31:0] p22_add_65458_comb;
  wire [31:0] p22_add_65480_comb;
  assign p22_and_65459_comb = p21_add_65377 & p21_add_65273;
  assign p22_add_65451_comb = (p21_add_65349 & p21_add_65248 ^ ~(p21_add_65349 | ~p21_add_65110)) + {p21_add_65349[5:0] ^ p21_add_65349[10:5] ^ p21_add_65349[24:19], p21_add_65349[31:27] ^ p21_add_65349[4:0] ^ p21_add_65349[18:14], p21_add_65349[26:13] ^ p21_add_65349[31:18] ^ p21_add_65349[13:0], p21_add_65349[12:6] ^ p21_add_65349[17:11] ^ p21_add_65349[31:25]};
  assign p22_add_65456_comb = p21_add_63845[31:2] + 30'h172c_2a77;
  assign p22_add_65452_comb = p22_add_65451_comb + p21_add_65355;
  assign p22_add_65478_comb = (p22_and_65459_comb ^ p21_add_65377 & p21_add_65137 ^ p21_and_65356) + p21_add_65348;
  assign p22_add_65453_comb = p22_add_65452_comb + p21_add_65137;
  assign p22_add_65458_comb = {p22_add_65456_comb, p21_bit_slice_64103} + p21_add_65110;
  assign p22_add_65480_comb = p22_add_65478_comb + {p21_add_65377[1:0] ^ p21_add_65377[12:11] ^ p21_add_65377[21:20], p21_add_65377[31:21] ^ p21_add_65377[10:0] ^ p21_add_65377[19:9], p21_add_65377[20:12] ^ p21_add_65377[31:23] ^ p21_add_65377[8:0], p21_add_65377[11:2] ^ p21_add_65377[22:13] ^ p21_add_65377[31:22]};

  // Registers for pipe stage 22:
  reg [31:0] p22_add_65248;
  reg [31:0] p22_add_63775;
  reg [31:0] p22_add_65349;
  reg [31:0] p22_add_64102;
  reg [31:0] p22_add_65452;
  reg [31:0] p22_add_65453;
  reg [31:0] p22_add_63845;
  reg [31:0] p22_add_65458;
  reg [31:0] p22_add_65273;
  reg [31:0] p22_add_64121;
  reg [31:0] p22_add_65377;
  reg [31:0] p22_add_64138;
  reg [31:0] p22_and_65459;
  reg [31:0] p22_add_65480;
  reg [31:0] p22_add_64290;
  reg [31:0] p22_add_64291;
  reg [31:0] p22_add_64441;
  reg [31:0] p22_add_64326;
  reg [31:0] p22_add_64459;
  reg [31:0] p22_add_64477;
  reg [31:0] p22_add_64612;
  reg [31:0] p22_add_64750;
  reg [31:0] p22_add_64891;
  reg [31:0] p22_add_65032;
  reg [31:0] p22_add_65172;
  always_ff @ (posedge clk) begin
    p22_add_65248 <= p21_add_65248;
    p22_add_63775 <= p21_add_63775;
    p22_add_65349 <= p21_add_65349;
    p22_add_64102 <= p21_add_64102;
    p22_add_65452 <= p22_add_65452_comb;
    p22_add_65453 <= p22_add_65453_comb;
    p22_add_63845 <= p21_add_63845;
    p22_add_65458 <= p22_add_65458_comb;
    p22_add_65273 <= p21_add_65273;
    p22_add_64121 <= p21_add_64121;
    p22_add_65377 <= p21_add_65377;
    p22_add_64138 <= p21_add_64138;
    p22_and_65459 <= p22_and_65459_comb;
    p22_add_65480 <= p22_add_65480_comb;
    p22_add_64290 <= p21_add_64290;
    p22_add_64291 <= p21_add_64291;
    p22_add_64441 <= p21_add_64441;
    p22_add_64326 <= p21_add_64326;
    p22_add_64459 <= p21_add_64459;
    p22_add_64477 <= p21_add_64477;
    p22_add_64612 <= p21_add_64612;
    p22_add_64750 <= p21_add_64750;
    p22_add_64891 <= p21_add_64891;
    p22_add_65032 <= p21_add_65032;
    p22_add_65172 <= p21_add_65172;
  end

  // ===== Pipe stage 23:
  wire [31:0] p23_and_65561_comb;
  wire [31:0] p23_add_65552_comb;
  wire [30:0] p23_add_65557_comb;
  wire [31:0] p23_add_65553_comb;
  wire [31:0] p23_add_65580_comb;
  wire [31:0] p23_add_65554_comb;
  wire [31:0] p23_add_65560_comb;
  wire [31:0] p23_add_65582_comb;
  assign p23_and_65561_comb = p22_add_65480 & p22_add_65377;
  assign p23_add_65552_comb = (p22_add_65453 & p22_add_65349 ^ ~(p22_add_65453 | ~p22_add_65248)) + {p22_add_65453[5:0] ^ p22_add_65453[10:5] ^ p22_add_65453[24:19], p22_add_65453[31:27] ^ p22_add_65453[4:0] ^ p22_add_65453[18:14], p22_add_65453[26:13] ^ p22_add_65453[31:18] ^ p22_add_65453[13:0], p22_add_65453[12:6] ^ p22_add_65453[17:11] ^ p22_add_65453[31:25]};
  assign p23_add_65557_comb = p22_add_64121[31:1] + 31'h3b7c_c46d;
  assign p23_add_65553_comb = p23_add_65552_comb + p22_add_65458;
  assign p23_add_65580_comb = (p23_and_65561_comb ^ p22_add_65480 & p22_add_65273 ^ p22_and_65459) + p22_add_65452;
  assign p23_add_65554_comb = p23_add_65553_comb + p22_add_65273;
  assign p23_add_65560_comb = {p23_add_65557_comb, p22_add_64121[0]} + p22_add_65248;
  assign p23_add_65582_comb = p23_add_65580_comb + {p22_add_65480[1:0] ^ p22_add_65480[12:11] ^ p22_add_65480[21:20], p22_add_65480[31:21] ^ p22_add_65480[10:0] ^ p22_add_65480[19:9], p22_add_65480[20:12] ^ p22_add_65480[31:23] ^ p22_add_65480[8:0], p22_add_65480[11:2] ^ p22_add_65480[22:13] ^ p22_add_65480[31:22]};

  // Registers for pipe stage 23:
  reg [31:0] p23_add_63775;
  reg [31:0] p23_add_65349;
  reg [31:0] p23_add_64102;
  reg [31:0] p23_add_65453;
  reg [31:0] p23_add_63845;
  reg [31:0] p23_add_65553;
  reg [31:0] p23_add_65554;
  reg [31:0] p23_add_64121;
  reg [31:0] p23_add_65560;
  reg [31:0] p23_add_65377;
  reg [31:0] p23_add_64138;
  reg [31:0] p23_add_65480;
  reg [31:0] p23_add_64290;
  reg [31:0] p23_and_65561;
  reg [31:0] p23_add_65582;
  reg [31:0] p23_add_64291;
  reg [31:0] p23_add_64441;
  reg [31:0] p23_add_64326;
  reg [31:0] p23_add_64459;
  reg [31:0] p23_add_64477;
  reg [31:0] p23_add_64612;
  reg [31:0] p23_add_64750;
  reg [31:0] p23_add_64891;
  reg [31:0] p23_add_65032;
  reg [31:0] p23_add_65172;
  always_ff @ (posedge clk) begin
    p23_add_63775 <= p22_add_63775;
    p23_add_65349 <= p22_add_65349;
    p23_add_64102 <= p22_add_64102;
    p23_add_65453 <= p22_add_65453;
    p23_add_63845 <= p22_add_63845;
    p23_add_65553 <= p23_add_65553_comb;
    p23_add_65554 <= p23_add_65554_comb;
    p23_add_64121 <= p22_add_64121;
    p23_add_65560 <= p23_add_65560_comb;
    p23_add_65377 <= p22_add_65377;
    p23_add_64138 <= p22_add_64138;
    p23_add_65480 <= p22_add_65480;
    p23_add_64290 <= p22_add_64290;
    p23_and_65561 <= p23_and_65561_comb;
    p23_add_65582 <= p23_add_65582_comb;
    p23_add_64291 <= p22_add_64291;
    p23_add_64441 <= p22_add_64441;
    p23_add_64326 <= p22_add_64326;
    p23_add_64459 <= p22_add_64459;
    p23_add_64477 <= p22_add_64477;
    p23_add_64612 <= p22_add_64612;
    p23_add_64750 <= p22_add_64750;
    p23_add_64891 <= p22_add_64891;
    p23_add_65032 <= p22_add_65032;
    p23_add_65172 <= p22_add_65172;
  end

  // ===== Pipe stage 24:
  wire [31:0] p24_and_65663_comb;
  wire [31:0] p24_add_65654_comb;
  wire [30:0] p24_add_65659_comb;
  wire [31:0] p24_add_65655_comb;
  wire [31:0] p24_add_65682_comb;
  wire [31:0] p24_add_65656_comb;
  wire [31:0] p24_add_65662_comb;
  wire [31:0] p24_add_65684_comb;
  assign p24_and_65663_comb = p23_add_65582 & p23_add_65480;
  assign p24_add_65654_comb = (p23_add_65554 & p23_add_65453 ^ ~(p23_add_65554 | ~p23_add_65349)) + {p23_add_65554[5:0] ^ p23_add_65554[10:5] ^ p23_add_65554[24:19], p23_add_65554[31:27] ^ p23_add_65554[4:0] ^ p23_add_65554[18:14], p23_add_65554[26:13] ^ p23_add_65554[31:18] ^ p23_add_65554[13:0], p23_add_65554[12:6] ^ p23_add_65554[17:11] ^ p23_add_65554[31:25]};
  assign p24_add_65659_comb = p23_add_64138[31:1] + 31'h4c1f_28a9;
  assign p24_add_65655_comb = p24_add_65654_comb + p23_add_65560;
  assign p24_add_65682_comb = (p24_and_65663_comb ^ p23_add_65582 & p23_add_65377 ^ p23_and_65561) + p23_add_65553;
  assign p24_add_65656_comb = p24_add_65655_comb + p23_add_65377;
  assign p24_add_65662_comb = {p24_add_65659_comb, p23_add_64138[0]} + p23_add_65349;
  assign p24_add_65684_comb = p24_add_65682_comb + {p23_add_65582[1:0] ^ p23_add_65582[12:11] ^ p23_add_65582[21:20], p23_add_65582[31:21] ^ p23_add_65582[10:0] ^ p23_add_65582[19:9], p23_add_65582[20:12] ^ p23_add_65582[31:23] ^ p23_add_65582[8:0], p23_add_65582[11:2] ^ p23_add_65582[22:13] ^ p23_add_65582[31:22]};

  // Registers for pipe stage 24:
  reg [31:0] p24_add_63775;
  reg [31:0] p24_add_64102;
  reg [31:0] p24_add_65453;
  reg [31:0] p24_add_63845;
  reg [31:0] p24_add_65554;
  reg [31:0] p24_add_64121;
  reg [31:0] p24_add_65655;
  reg [31:0] p24_add_65656;
  reg [31:0] p24_add_64138;
  reg [31:0] p24_add_65662;
  reg [31:0] p24_add_65480;
  reg [31:0] p24_add_64290;
  reg [31:0] p24_add_65582;
  reg [31:0] p24_add_64291;
  reg [31:0] p24_and_65663;
  reg [31:0] p24_add_65684;
  reg [31:0] p24_add_64441;
  reg [31:0] p24_add_64326;
  reg [31:0] p24_add_64459;
  reg [31:0] p24_add_64477;
  reg [31:0] p24_add_64612;
  reg [31:0] p24_add_64750;
  reg [31:0] p24_add_64891;
  reg [31:0] p24_add_65032;
  reg [31:0] p24_add_65172;
  always_ff @ (posedge clk) begin
    p24_add_63775 <= p23_add_63775;
    p24_add_64102 <= p23_add_64102;
    p24_add_65453 <= p23_add_65453;
    p24_add_63845 <= p23_add_63845;
    p24_add_65554 <= p23_add_65554;
    p24_add_64121 <= p23_add_64121;
    p24_add_65655 <= p24_add_65655_comb;
    p24_add_65656 <= p24_add_65656_comb;
    p24_add_64138 <= p23_add_64138;
    p24_add_65662 <= p24_add_65662_comb;
    p24_add_65480 <= p23_add_65480;
    p24_add_64290 <= p23_add_64290;
    p24_add_65582 <= p23_add_65582;
    p24_add_64291 <= p23_add_64291;
    p24_and_65663 <= p24_and_65663_comb;
    p24_add_65684 <= p24_add_65684_comb;
    p24_add_64441 <= p23_add_64441;
    p24_add_64326 <= p23_add_64326;
    p24_add_64459 <= p23_add_64459;
    p24_add_64477 <= p23_add_64477;
    p24_add_64612 <= p23_add_64612;
    p24_add_64750 <= p23_add_64750;
    p24_add_64891 <= p23_add_64891;
    p24_add_65032 <= p23_add_65032;
    p24_add_65172 <= p23_add_65172;
  end

  // ===== Pipe stage 25:
  wire [31:0] p25_and_65762_comb;
  wire [31:0] p25_add_65756_comb;
  wire [31:0] p25_add_65757_comb;
  wire [31:0] p25_add_65760_comb;
  wire [31:0] p25_add_65781_comb;
  wire [31:0] p25_add_65758_comb;
  wire [31:0] p25_add_65761_comb;
  wire [31:0] p25_add_65783_comb;
  assign p25_and_65762_comb = p24_add_65684 & p24_add_65582;
  assign p25_add_65756_comb = (p24_add_65656 & p24_add_65554 ^ ~(p24_add_65656 | ~p24_add_65453)) + {p24_add_65656[5:0] ^ p24_add_65656[10:5] ^ p24_add_65656[24:19], p24_add_65656[31:27] ^ p24_add_65656[4:0] ^ p24_add_65656[18:14], p24_add_65656[26:13] ^ p24_add_65656[31:18] ^ p24_add_65656[13:0], p24_add_65656[12:6] ^ p24_add_65656[17:11] ^ p24_add_65656[31:25]};
  assign p25_add_65757_comb = p25_add_65756_comb + p24_add_65662;
  assign p25_add_65760_comb = p24_add_64290 + 32'ha831_c66d;
  assign p25_add_65781_comb = (p25_and_65762_comb ^ p24_add_65684 & p24_add_65480 ^ p24_and_65663) + p24_add_65655;
  assign p25_add_65758_comb = p25_add_65757_comb + p24_add_65480;
  assign p25_add_65761_comb = p24_add_65453 + p25_add_65760_comb;
  assign p25_add_65783_comb = p25_add_65781_comb + {p24_add_65684[1:0] ^ p24_add_65684[12:11] ^ p24_add_65684[21:20], p24_add_65684[31:21] ^ p24_add_65684[10:0] ^ p24_add_65684[19:9], p24_add_65684[20:12] ^ p24_add_65684[31:23] ^ p24_add_65684[8:0], p24_add_65684[11:2] ^ p24_add_65684[22:13] ^ p24_add_65684[31:22]};

  // Registers for pipe stage 25:
  reg [31:0] p25_add_63775;
  reg [31:0] p25_add_64102;
  reg [31:0] p25_add_63845;
  reg [31:0] p25_add_65554;
  reg [31:0] p25_add_64121;
  reg [31:0] p25_add_65656;
  reg [31:0] p25_add_64138;
  reg [31:0] p25_add_65757;
  reg [31:0] p25_add_65758;
  reg [31:0] p25_add_64290;
  reg [31:0] p25_add_65761;
  reg [31:0] p25_add_65582;
  reg [31:0] p25_add_64291;
  reg [31:0] p25_add_65684;
  reg [31:0] p25_add_64441;
  reg [31:0] p25_and_65762;
  reg [31:0] p25_add_65783;
  reg [31:0] p25_add_64326;
  reg [31:0] p25_add_64459;
  reg [31:0] p25_add_64477;
  reg [31:0] p25_add_64612;
  reg [31:0] p25_add_64750;
  reg [31:0] p25_add_64891;
  reg [31:0] p25_add_65032;
  reg [31:0] p25_add_65172;
  always_ff @ (posedge clk) begin
    p25_add_63775 <= p24_add_63775;
    p25_add_64102 <= p24_add_64102;
    p25_add_63845 <= p24_add_63845;
    p25_add_65554 <= p24_add_65554;
    p25_add_64121 <= p24_add_64121;
    p25_add_65656 <= p24_add_65656;
    p25_add_64138 <= p24_add_64138;
    p25_add_65757 <= p25_add_65757_comb;
    p25_add_65758 <= p25_add_65758_comb;
    p25_add_64290 <= p24_add_64290;
    p25_add_65761 <= p25_add_65761_comb;
    p25_add_65582 <= p24_add_65582;
    p25_add_64291 <= p24_add_64291;
    p25_add_65684 <= p24_add_65684;
    p25_add_64441 <= p24_add_64441;
    p25_and_65762 <= p25_and_65762_comb;
    p25_add_65783 <= p25_add_65783_comb;
    p25_add_64326 <= p24_add_64326;
    p25_add_64459 <= p24_add_64459;
    p25_add_64477 <= p24_add_64477;
    p25_add_64612 <= p24_add_64612;
    p25_add_64750 <= p24_add_64750;
    p25_add_64891 <= p24_add_64891;
    p25_add_65032 <= p24_add_65032;
    p25_add_65172 <= p24_add_65172;
  end

  // ===== Pipe stage 26:
  wire [31:0] p26_and_65864_comb;
  wire [31:0] p26_add_65855_comb;
  wire [28:0] p26_add_65860_comb;
  wire [31:0] p26_add_65856_comb;
  wire [31:0] p26_add_65883_comb;
  wire [31:0] p26_add_65857_comb;
  wire [31:0] p26_add_65863_comb;
  wire [31:0] p26_add_65885_comb;
  assign p26_and_65864_comb = p25_add_65783 & p25_add_65684;
  assign p26_add_65855_comb = {p25_add_65758[5:0] ^ p25_add_65758[10:5] ^ p25_add_65758[24:19], p25_add_65758[31:27] ^ p25_add_65758[4:0] ^ p25_add_65758[18:14], p25_add_65758[26:13] ^ p25_add_65758[31:18] ^ p25_add_65758[13:0], p25_add_65758[12:6] ^ p25_add_65758[17:11] ^ p25_add_65758[31:25]} + (p25_add_65758 & p25_add_65656 ^ ~(p25_add_65758 | ~p25_add_65554));
  assign p26_add_65860_comb = p25_add_64291[31:3] + 29'h1600_64f9;
  assign p26_add_65856_comb = p26_add_65855_comb + p25_add_65761;
  assign p26_add_65883_comb = (p26_and_65864_comb ^ p25_add_65783 & p25_add_65582 ^ p25_and_65762) + p25_add_65757;
  assign p26_add_65857_comb = p26_add_65856_comb + p25_add_65582;
  assign p26_add_65863_comb = {p26_add_65860_comb, p25_add_64291[2:0]} + p25_add_65554;
  assign p26_add_65885_comb = p26_add_65883_comb + {p25_add_65783[1:0] ^ p25_add_65783[12:11] ^ p25_add_65783[21:20], p25_add_65783[31:21] ^ p25_add_65783[10:0] ^ p25_add_65783[19:9], p25_add_65783[20:12] ^ p25_add_65783[31:23] ^ p25_add_65783[8:0], p25_add_65783[11:2] ^ p25_add_65783[22:13] ^ p25_add_65783[31:22]};

  // Registers for pipe stage 26:
  reg [31:0] p26_add_63775;
  reg [31:0] p26_add_64102;
  reg [31:0] p26_add_63845;
  reg [31:0] p26_add_64121;
  reg [31:0] p26_add_65656;
  reg [31:0] p26_add_64138;
  reg [31:0] p26_add_65758;
  reg [31:0] p26_add_64290;
  reg [31:0] p26_add_65856;
  reg [31:0] p26_add_65857;
  reg [31:0] p26_add_64291;
  reg [31:0] p26_add_65863;
  reg [31:0] p26_add_65684;
  reg [31:0] p26_add_64441;
  reg [31:0] p26_add_65783;
  reg [31:0] p26_add_64326;
  reg [31:0] p26_and_65864;
  reg [31:0] p26_add_65885;
  reg [31:0] p26_add_64459;
  reg [31:0] p26_add_64477;
  reg [31:0] p26_add_64612;
  reg [31:0] p26_add_64750;
  reg [31:0] p26_add_64891;
  reg [31:0] p26_add_65032;
  reg [31:0] p26_add_65172;
  always_ff @ (posedge clk) begin
    p26_add_63775 <= p25_add_63775;
    p26_add_64102 <= p25_add_64102;
    p26_add_63845 <= p25_add_63845;
    p26_add_64121 <= p25_add_64121;
    p26_add_65656 <= p25_add_65656;
    p26_add_64138 <= p25_add_64138;
    p26_add_65758 <= p25_add_65758;
    p26_add_64290 <= p25_add_64290;
    p26_add_65856 <= p26_add_65856_comb;
    p26_add_65857 <= p26_add_65857_comb;
    p26_add_64291 <= p25_add_64291;
    p26_add_65863 <= p26_add_65863_comb;
    p26_add_65684 <= p25_add_65684;
    p26_add_64441 <= p25_add_64441;
    p26_add_65783 <= p25_add_65783;
    p26_add_64326 <= p25_add_64326;
    p26_and_65864 <= p26_and_65864_comb;
    p26_add_65885 <= p26_add_65885_comb;
    p26_add_64459 <= p25_add_64459;
    p26_add_64477 <= p25_add_64477;
    p26_add_64612 <= p25_add_64612;
    p26_add_64750 <= p25_add_64750;
    p26_add_64891 <= p25_add_64891;
    p26_add_65032 <= p25_add_65032;
    p26_add_65172 <= p25_add_65172;
  end

  // ===== Pipe stage 27:
  wire [31:0] p27_and_65963_comb;
  wire [31:0] p27_add_65957_comb;
  wire [31:0] p27_add_65958_comb;
  wire [31:0] p27_add_65961_comb;
  wire [31:0] p27_add_65982_comb;
  wire [31:0] p27_add_65959_comb;
  wire [31:0] p27_add_65962_comb;
  wire [31:0] p27_add_65984_comb;
  assign p27_and_65963_comb = p26_add_65885 & p26_add_65783;
  assign p27_add_65957_comb = (p26_add_65857 & p26_add_65758 ^ ~(p26_add_65857 | ~p26_add_65656)) + {p26_add_65857[5:0] ^ p26_add_65857[10:5] ^ p26_add_65857[24:19], p26_add_65857[31:27] ^ p26_add_65857[4:0] ^ p26_add_65857[18:14], p26_add_65857[26:13] ^ p26_add_65857[31:18] ^ p26_add_65857[13:0], p26_add_65857[12:6] ^ p26_add_65857[17:11] ^ p26_add_65857[31:25]};
  assign p27_add_65958_comb = p27_add_65957_comb + p26_add_65863;
  assign p27_add_65961_comb = p26_add_64441 + 32'hbf59_7fc7;
  assign p27_add_65982_comb = (p27_and_65963_comb ^ p26_add_65885 & p26_add_65684 ^ p26_and_65864) + p26_add_65856;
  assign p27_add_65959_comb = p27_add_65958_comb + p26_add_65684;
  assign p27_add_65962_comb = p26_add_65656 + p27_add_65961_comb;
  assign p27_add_65984_comb = p27_add_65982_comb + {p26_add_65885[1:0] ^ p26_add_65885[12:11] ^ p26_add_65885[21:20], p26_add_65885[31:21] ^ p26_add_65885[10:0] ^ p26_add_65885[19:9], p26_add_65885[20:12] ^ p26_add_65885[31:23] ^ p26_add_65885[8:0], p26_add_65885[11:2] ^ p26_add_65885[22:13] ^ p26_add_65885[31:22]};

  // Registers for pipe stage 27:
  reg [31:0] p27_add_63775;
  reg [31:0] p27_add_64102;
  reg [31:0] p27_add_63845;
  reg [31:0] p27_add_64121;
  reg [31:0] p27_add_64138;
  reg [31:0] p27_add_65758;
  reg [31:0] p27_add_64290;
  reg [31:0] p27_add_65857;
  reg [31:0] p27_add_64291;
  reg [31:0] p27_add_65958;
  reg [31:0] p27_add_65959;
  reg [31:0] p27_add_64441;
  reg [31:0] p27_add_65962;
  reg [31:0] p27_add_65783;
  reg [31:0] p27_add_64326;
  reg [31:0] p27_add_65885;
  reg [31:0] p27_add_64459;
  reg [31:0] p27_and_65963;
  reg [31:0] p27_add_65984;
  reg [31:0] p27_add_64477;
  reg [31:0] p27_add_64612;
  reg [31:0] p27_add_64750;
  reg [31:0] p27_add_64891;
  reg [31:0] p27_add_65032;
  reg [31:0] p27_add_65172;
  always_ff @ (posedge clk) begin
    p27_add_63775 <= p26_add_63775;
    p27_add_64102 <= p26_add_64102;
    p27_add_63845 <= p26_add_63845;
    p27_add_64121 <= p26_add_64121;
    p27_add_64138 <= p26_add_64138;
    p27_add_65758 <= p26_add_65758;
    p27_add_64290 <= p26_add_64290;
    p27_add_65857 <= p26_add_65857;
    p27_add_64291 <= p26_add_64291;
    p27_add_65958 <= p27_add_65958_comb;
    p27_add_65959 <= p27_add_65959_comb;
    p27_add_64441 <= p26_add_64441;
    p27_add_65962 <= p27_add_65962_comb;
    p27_add_65783 <= p26_add_65783;
    p27_add_64326 <= p26_add_64326;
    p27_add_65885 <= p26_add_65885;
    p27_add_64459 <= p26_add_64459;
    p27_and_65963 <= p27_and_65963_comb;
    p27_add_65984 <= p27_add_65984_comb;
    p27_add_64477 <= p26_add_64477;
    p27_add_64612 <= p26_add_64612;
    p27_add_64750 <= p26_add_64750;
    p27_add_64891 <= p26_add_64891;
    p27_add_65032 <= p26_add_65032;
    p27_add_65172 <= p26_add_65172;
  end

  // ===== Pipe stage 28:
  wire [31:0] p28_and_66062_comb;
  wire [31:0] p28_add_66056_comb;
  wire [31:0] p28_add_66057_comb;
  wire [31:0] p28_add_66060_comb;
  wire [31:0] p28_add_66081_comb;
  wire [31:0] p28_add_66058_comb;
  wire [31:0] p28_add_66061_comb;
  wire [31:0] p28_add_66083_comb;
  assign p28_and_66062_comb = p27_add_65984 & p27_add_65885;
  assign p28_add_66056_comb = {p27_add_65959[5:0] ^ p27_add_65959[10:5] ^ p27_add_65959[24:19], p27_add_65959[31:27] ^ p27_add_65959[4:0] ^ p27_add_65959[18:14], p27_add_65959[26:13] ^ p27_add_65959[31:18] ^ p27_add_65959[13:0], p27_add_65959[12:6] ^ p27_add_65959[17:11] ^ p27_add_65959[31:25]} + (p27_add_65959 & p27_add_65857 ^ ~(p27_add_65959 | ~p27_add_65758));
  assign p28_add_66057_comb = p28_add_66056_comb + p27_add_65962;
  assign p28_add_66060_comb = p27_add_64326 + 32'hc6e0_0bf3;
  assign p28_add_66081_comb = (p28_and_66062_comb ^ p27_add_65984 & p27_add_65783 ^ p27_and_65963) + p27_add_65958;
  assign p28_add_66058_comb = p28_add_66057_comb + p27_add_65783;
  assign p28_add_66061_comb = p27_add_65758 + p28_add_66060_comb;
  assign p28_add_66083_comb = p28_add_66081_comb + {p27_add_65984[1:0] ^ p27_add_65984[12:11] ^ p27_add_65984[21:20], p27_add_65984[31:21] ^ p27_add_65984[10:0] ^ p27_add_65984[19:9], p27_add_65984[20:12] ^ p27_add_65984[31:23] ^ p27_add_65984[8:0], p27_add_65984[11:2] ^ p27_add_65984[22:13] ^ p27_add_65984[31:22]};

  // Registers for pipe stage 28:
  reg [31:0] p28_add_63775;
  reg [31:0] p28_add_64102;
  reg [31:0] p28_add_63845;
  reg [31:0] p28_add_64121;
  reg [31:0] p28_add_64138;
  reg [31:0] p28_add_64290;
  reg [31:0] p28_add_65857;
  reg [31:0] p28_add_64291;
  reg [31:0] p28_add_65959;
  reg [31:0] p28_add_64441;
  reg [31:0] p28_add_66057;
  reg [31:0] p28_add_66058;
  reg [31:0] p28_add_64326;
  reg [31:0] p28_add_66061;
  reg [31:0] p28_add_65885;
  reg [31:0] p28_add_64459;
  reg [31:0] p28_add_65984;
  reg [31:0] p28_add_64477;
  reg [31:0] p28_and_66062;
  reg [31:0] p28_add_66083;
  reg [31:0] p28_add_64612;
  reg [31:0] p28_add_64750;
  reg [31:0] p28_add_64891;
  reg [31:0] p28_add_65032;
  reg [31:0] p28_add_65172;
  always_ff @ (posedge clk) begin
    p28_add_63775 <= p27_add_63775;
    p28_add_64102 <= p27_add_64102;
    p28_add_63845 <= p27_add_63845;
    p28_add_64121 <= p27_add_64121;
    p28_add_64138 <= p27_add_64138;
    p28_add_64290 <= p27_add_64290;
    p28_add_65857 <= p27_add_65857;
    p28_add_64291 <= p27_add_64291;
    p28_add_65959 <= p27_add_65959;
    p28_add_64441 <= p27_add_64441;
    p28_add_66057 <= p28_add_66057_comb;
    p28_add_66058 <= p28_add_66058_comb;
    p28_add_64326 <= p27_add_64326;
    p28_add_66061 <= p28_add_66061_comb;
    p28_add_65885 <= p27_add_65885;
    p28_add_64459 <= p27_add_64459;
    p28_add_65984 <= p27_add_65984;
    p28_add_64477 <= p27_add_64477;
    p28_and_66062 <= p28_and_66062_comb;
    p28_add_66083 <= p28_add_66083_comb;
    p28_add_64612 <= p27_add_64612;
    p28_add_64750 <= p27_add_64750;
    p28_add_64891 <= p27_add_64891;
    p28_add_65032 <= p27_add_65032;
    p28_add_65172 <= p27_add_65172;
  end

  // ===== Pipe stage 29:
  wire [31:0] p29_and_66161_comb;
  wire [31:0] p29_add_66155_comb;
  wire [31:0] p29_add_66156_comb;
  wire [31:0] p29_add_66159_comb;
  wire [31:0] p29_add_66180_comb;
  wire [31:0] p29_add_66157_comb;
  wire [31:0] p29_add_66160_comb;
  wire [31:0] p29_add_66182_comb;
  assign p29_and_66161_comb = p28_add_66083 & p28_add_65984;
  assign p29_add_66155_comb = {p28_add_66058[5:0] ^ p28_add_66058[10:5] ^ p28_add_66058[24:19], p28_add_66058[31:27] ^ p28_add_66058[4:0] ^ p28_add_66058[18:14], p28_add_66058[26:13] ^ p28_add_66058[31:18] ^ p28_add_66058[13:0], p28_add_66058[12:6] ^ p28_add_66058[17:11] ^ p28_add_66058[31:25]} + (p28_add_66058 & p28_add_65959 ^ ~(p28_add_66058 | ~p28_add_65857));
  assign p29_add_66156_comb = p29_add_66155_comb + p28_add_66061;
  assign p29_add_66159_comb = p28_add_64459 + 32'hd5a7_9147;
  assign p29_add_66180_comb = (p29_and_66161_comb ^ p28_add_66083 & p28_add_65885 ^ p28_and_66062) + p28_add_66057;
  assign p29_add_66157_comb = p29_add_66156_comb + p28_add_65885;
  assign p29_add_66160_comb = p28_add_65857 + p29_add_66159_comb;
  assign p29_add_66182_comb = p29_add_66180_comb + {p28_add_66083[1:0] ^ p28_add_66083[12:11] ^ p28_add_66083[21:20], p28_add_66083[31:21] ^ p28_add_66083[10:0] ^ p28_add_66083[19:9], p28_add_66083[20:12] ^ p28_add_66083[31:23] ^ p28_add_66083[8:0], p28_add_66083[11:2] ^ p28_add_66083[22:13] ^ p28_add_66083[31:22]};

  // Registers for pipe stage 29:
  reg [31:0] p29_add_63775;
  reg [31:0] p29_add_64102;
  reg [31:0] p29_add_63845;
  reg [31:0] p29_add_64121;
  reg [31:0] p29_add_64138;
  reg [31:0] p29_add_64290;
  reg [31:0] p29_add_64291;
  reg [31:0] p29_add_65959;
  reg [31:0] p29_add_64441;
  reg [31:0] p29_add_66058;
  reg [31:0] p29_add_64326;
  reg [31:0] p29_add_66156;
  reg [31:0] p29_add_66157;
  reg [31:0] p29_add_64459;
  reg [31:0] p29_add_66160;
  reg [31:0] p29_add_65984;
  reg [31:0] p29_add_64477;
  reg [31:0] p29_add_66083;
  reg [31:0] p29_add_64612;
  reg [31:0] p29_and_66161;
  reg [31:0] p29_add_66182;
  reg [31:0] p29_add_64750;
  reg [31:0] p29_add_64891;
  reg [31:0] p29_add_65032;
  reg [31:0] p29_add_65172;
  always_ff @ (posedge clk) begin
    p29_add_63775 <= p28_add_63775;
    p29_add_64102 <= p28_add_64102;
    p29_add_63845 <= p28_add_63845;
    p29_add_64121 <= p28_add_64121;
    p29_add_64138 <= p28_add_64138;
    p29_add_64290 <= p28_add_64290;
    p29_add_64291 <= p28_add_64291;
    p29_add_65959 <= p28_add_65959;
    p29_add_64441 <= p28_add_64441;
    p29_add_66058 <= p28_add_66058;
    p29_add_64326 <= p28_add_64326;
    p29_add_66156 <= p29_add_66156_comb;
    p29_add_66157 <= p29_add_66157_comb;
    p29_add_64459 <= p28_add_64459;
    p29_add_66160 <= p29_add_66160_comb;
    p29_add_65984 <= p28_add_65984;
    p29_add_64477 <= p28_add_64477;
    p29_add_66083 <= p28_add_66083;
    p29_add_64612 <= p28_add_64612;
    p29_and_66161 <= p29_and_66161_comb;
    p29_add_66182 <= p29_add_66182_comb;
    p29_add_64750 <= p28_add_64750;
    p29_add_64891 <= p28_add_64891;
    p29_add_65032 <= p28_add_65032;
    p29_add_65172 <= p28_add_65172;
  end

  // ===== Pipe stage 30:
  wire [31:0] p30_and_66260_comb;
  wire [31:0] p30_add_66254_comb;
  wire [31:0] p30_add_66255_comb;
  wire [31:0] p30_add_66258_comb;
  wire [31:0] p30_add_66279_comb;
  wire [31:0] p30_add_66256_comb;
  wire [31:0] p30_add_66259_comb;
  wire [31:0] p30_add_66281_comb;
  assign p30_and_66260_comb = p29_add_66182 & p29_add_66083;
  assign p30_add_66254_comb = {p29_add_66157[5:0] ^ p29_add_66157[10:5] ^ p29_add_66157[24:19], p29_add_66157[31:27] ^ p29_add_66157[4:0] ^ p29_add_66157[18:14], p29_add_66157[26:13] ^ p29_add_66157[31:18] ^ p29_add_66157[13:0], p29_add_66157[12:6] ^ p29_add_66157[17:11] ^ p29_add_66157[31:25]} + (p29_add_66157 & p29_add_66058 ^ ~(p29_add_66157 | ~p29_add_65959));
  assign p30_add_66255_comb = p30_add_66254_comb + p29_add_66160;
  assign p30_add_66258_comb = p29_add_64477 + 32'h06ca_6351;
  assign p30_add_66279_comb = (p30_and_66260_comb ^ p29_add_66182 & p29_add_65984 ^ p29_and_66161) + p29_add_66156;
  assign p30_add_66256_comb = p30_add_66255_comb + p29_add_65984;
  assign p30_add_66259_comb = p29_add_65959 + p30_add_66258_comb;
  assign p30_add_66281_comb = p30_add_66279_comb + {p29_add_66182[1:0] ^ p29_add_66182[12:11] ^ p29_add_66182[21:20], p29_add_66182[31:21] ^ p29_add_66182[10:0] ^ p29_add_66182[19:9], p29_add_66182[20:12] ^ p29_add_66182[31:23] ^ p29_add_66182[8:0], p29_add_66182[11:2] ^ p29_add_66182[22:13] ^ p29_add_66182[31:22]};

  // Registers for pipe stage 30:
  reg [31:0] p30_add_63775;
  reg [31:0] p30_add_64102;
  reg [31:0] p30_add_63845;
  reg [31:0] p30_add_64121;
  reg [31:0] p30_add_64138;
  reg [31:0] p30_add_64290;
  reg [31:0] p30_add_64291;
  reg [31:0] p30_add_64441;
  reg [31:0] p30_add_66058;
  reg [31:0] p30_add_64326;
  reg [31:0] p30_add_66157;
  reg [31:0] p30_add_64459;
  reg [31:0] p30_add_66255;
  reg [31:0] p30_add_66256;
  reg [31:0] p30_add_64477;
  reg [31:0] p30_add_66259;
  reg [31:0] p30_add_66083;
  reg [31:0] p30_add_64612;
  reg [31:0] p30_add_66182;
  reg [31:0] p30_add_64750;
  reg [31:0] p30_and_66260;
  reg [31:0] p30_add_66281;
  reg [31:0] p30_add_64891;
  reg [31:0] p30_add_65032;
  reg [31:0] p30_add_65172;
  always_ff @ (posedge clk) begin
    p30_add_63775 <= p29_add_63775;
    p30_add_64102 <= p29_add_64102;
    p30_add_63845 <= p29_add_63845;
    p30_add_64121 <= p29_add_64121;
    p30_add_64138 <= p29_add_64138;
    p30_add_64290 <= p29_add_64290;
    p30_add_64291 <= p29_add_64291;
    p30_add_64441 <= p29_add_64441;
    p30_add_66058 <= p29_add_66058;
    p30_add_64326 <= p29_add_64326;
    p30_add_66157 <= p29_add_66157;
    p30_add_64459 <= p29_add_64459;
    p30_add_66255 <= p30_add_66255_comb;
    p30_add_66256 <= p30_add_66256_comb;
    p30_add_64477 <= p29_add_64477;
    p30_add_66259 <= p30_add_66259_comb;
    p30_add_66083 <= p29_add_66083;
    p30_add_64612 <= p29_add_64612;
    p30_add_66182 <= p29_add_66182;
    p30_add_64750 <= p29_add_64750;
    p30_and_66260 <= p30_and_66260_comb;
    p30_add_66281 <= p30_add_66281_comb;
    p30_add_64891 <= p29_add_64891;
    p30_add_65032 <= p29_add_65032;
    p30_add_65172 <= p29_add_65172;
  end

  // ===== Pipe stage 31:
  wire [31:0] p31_and_66359_comb;
  wire [31:0] p31_add_66353_comb;
  wire [31:0] p31_add_66354_comb;
  wire [31:0] p31_add_66357_comb;
  wire [31:0] p31_add_66378_comb;
  wire [31:0] p31_add_66355_comb;
  wire [31:0] p31_add_66358_comb;
  wire [31:0] p31_add_66380_comb;
  assign p31_and_66359_comb = p30_add_66281 & p30_add_66182;
  assign p31_add_66353_comb = {p30_add_66256[5:0] ^ p30_add_66256[10:5] ^ p30_add_66256[24:19], p30_add_66256[31:27] ^ p30_add_66256[4:0] ^ p30_add_66256[18:14], p30_add_66256[26:13] ^ p30_add_66256[31:18] ^ p30_add_66256[13:0], p30_add_66256[12:6] ^ p30_add_66256[17:11] ^ p30_add_66256[31:25]} + (p30_add_66256 & p30_add_66157 ^ ~(p30_add_66256 | ~p30_add_66058));
  assign p31_add_66354_comb = p31_add_66353_comb + p30_add_66259;
  assign p31_add_66357_comb = p30_add_64612 + 32'h1429_2967;
  assign p31_add_66378_comb = (p31_and_66359_comb ^ p30_add_66281 & p30_add_66083 ^ p30_and_66260) + p30_add_66255;
  assign p31_add_66355_comb = p31_add_66354_comb + p30_add_66083;
  assign p31_add_66358_comb = p30_add_66058 + p31_add_66357_comb;
  assign p31_add_66380_comb = p31_add_66378_comb + {p30_add_66281[1:0] ^ p30_add_66281[12:11] ^ p30_add_66281[21:20], p30_add_66281[31:21] ^ p30_add_66281[10:0] ^ p30_add_66281[19:9], p30_add_66281[20:12] ^ p30_add_66281[31:23] ^ p30_add_66281[8:0], p30_add_66281[11:2] ^ p30_add_66281[22:13] ^ p30_add_66281[31:22]};

  // Registers for pipe stage 31:
  reg [31:0] p31_add_63775;
  reg [31:0] p31_add_64102;
  reg [31:0] p31_add_63845;
  reg [31:0] p31_add_64121;
  reg [31:0] p31_add_64138;
  reg [31:0] p31_add_64290;
  reg [31:0] p31_add_64291;
  reg [31:0] p31_add_64441;
  reg [31:0] p31_add_64326;
  reg [31:0] p31_add_66157;
  reg [31:0] p31_add_64459;
  reg [31:0] p31_add_66256;
  reg [31:0] p31_add_64477;
  reg [31:0] p31_add_66354;
  reg [31:0] p31_add_66355;
  reg [31:0] p31_add_64612;
  reg [31:0] p31_add_66358;
  reg [31:0] p31_add_66182;
  reg [31:0] p31_add_64750;
  reg [31:0] p31_add_66281;
  reg [31:0] p31_add_64891;
  reg [31:0] p31_and_66359;
  reg [31:0] p31_add_66380;
  reg [31:0] p31_add_65032;
  reg [31:0] p31_add_65172;
  always_ff @ (posedge clk) begin
    p31_add_63775 <= p30_add_63775;
    p31_add_64102 <= p30_add_64102;
    p31_add_63845 <= p30_add_63845;
    p31_add_64121 <= p30_add_64121;
    p31_add_64138 <= p30_add_64138;
    p31_add_64290 <= p30_add_64290;
    p31_add_64291 <= p30_add_64291;
    p31_add_64441 <= p30_add_64441;
    p31_add_64326 <= p30_add_64326;
    p31_add_66157 <= p30_add_66157;
    p31_add_64459 <= p30_add_64459;
    p31_add_66256 <= p30_add_66256;
    p31_add_64477 <= p30_add_64477;
    p31_add_66354 <= p31_add_66354_comb;
    p31_add_66355 <= p31_add_66355_comb;
    p31_add_64612 <= p30_add_64612;
    p31_add_66358 <= p31_add_66358_comb;
    p31_add_66182 <= p30_add_66182;
    p31_add_64750 <= p30_add_64750;
    p31_add_66281 <= p30_add_66281;
    p31_add_64891 <= p30_add_64891;
    p31_and_66359 <= p31_and_66359_comb;
    p31_add_66380 <= p31_add_66380_comb;
    p31_add_65032 <= p30_add_65032;
    p31_add_65172 <= p30_add_65172;
  end

  // ===== Pipe stage 32:
  wire [31:0] p32_and_66458_comb;
  wire [31:0] p32_add_66452_comb;
  wire [31:0] p32_add_66453_comb;
  wire [31:0] p32_add_66456_comb;
  wire [31:0] p32_add_66477_comb;
  wire [31:0] p32_add_66454_comb;
  wire [31:0] p32_add_66457_comb;
  wire [31:0] p32_add_66479_comb;
  assign p32_and_66458_comb = p31_add_66380 & p31_add_66281;
  assign p32_add_66452_comb = {p31_add_66355[5:0] ^ p31_add_66355[10:5] ^ p31_add_66355[24:19], p31_add_66355[31:27] ^ p31_add_66355[4:0] ^ p31_add_66355[18:14], p31_add_66355[26:13] ^ p31_add_66355[31:18] ^ p31_add_66355[13:0], p31_add_66355[12:6] ^ p31_add_66355[17:11] ^ p31_add_66355[31:25]} + (p31_add_66355 & p31_add_66256 ^ ~(p31_add_66355 | ~p31_add_66157));
  assign p32_add_66453_comb = p32_add_66452_comb + p31_add_66358;
  assign p32_add_66456_comb = p31_add_64750 + 32'h27b7_0a85;
  assign p32_add_66477_comb = (p32_and_66458_comb ^ p31_add_66380 & p31_add_66182 ^ p31_and_66359) + p31_add_66354;
  assign p32_add_66454_comb = p32_add_66453_comb + p31_add_66182;
  assign p32_add_66457_comb = p31_add_66157 + p32_add_66456_comb;
  assign p32_add_66479_comb = p32_add_66477_comb + {p31_add_66380[1:0] ^ p31_add_66380[12:11] ^ p31_add_66380[21:20], p31_add_66380[31:21] ^ p31_add_66380[10:0] ^ p31_add_66380[19:9], p31_add_66380[20:12] ^ p31_add_66380[31:23] ^ p31_add_66380[8:0], p31_add_66380[11:2] ^ p31_add_66380[22:13] ^ p31_add_66380[31:22]};

  // Registers for pipe stage 32:
  reg [31:0] p32_add_63775;
  reg [31:0] p32_add_64102;
  reg [31:0] p32_add_63845;
  reg [31:0] p32_add_64121;
  reg [31:0] p32_add_64138;
  reg [31:0] p32_add_64290;
  reg [31:0] p32_add_64291;
  reg [31:0] p32_add_64441;
  reg [31:0] p32_add_64326;
  reg [31:0] p32_add_64459;
  reg [31:0] p32_add_66256;
  reg [31:0] p32_add_64477;
  reg [31:0] p32_add_66355;
  reg [31:0] p32_add_64612;
  reg [31:0] p32_add_66453;
  reg [31:0] p32_add_66454;
  reg [31:0] p32_add_64750;
  reg [31:0] p32_add_66457;
  reg [31:0] p32_add_66281;
  reg [31:0] p32_add_64891;
  reg [31:0] p32_add_66380;
  reg [31:0] p32_add_65032;
  reg [31:0] p32_and_66458;
  reg [31:0] p32_add_66479;
  reg [31:0] p32_add_65172;
  always_ff @ (posedge clk) begin
    p32_add_63775 <= p31_add_63775;
    p32_add_64102 <= p31_add_64102;
    p32_add_63845 <= p31_add_63845;
    p32_add_64121 <= p31_add_64121;
    p32_add_64138 <= p31_add_64138;
    p32_add_64290 <= p31_add_64290;
    p32_add_64291 <= p31_add_64291;
    p32_add_64441 <= p31_add_64441;
    p32_add_64326 <= p31_add_64326;
    p32_add_64459 <= p31_add_64459;
    p32_add_66256 <= p31_add_66256;
    p32_add_64477 <= p31_add_64477;
    p32_add_66355 <= p31_add_66355;
    p32_add_64612 <= p31_add_64612;
    p32_add_66453 <= p32_add_66453_comb;
    p32_add_66454 <= p32_add_66454_comb;
    p32_add_64750 <= p31_add_64750;
    p32_add_66457 <= p32_add_66457_comb;
    p32_add_66281 <= p31_add_66281;
    p32_add_64891 <= p31_add_64891;
    p32_add_66380 <= p31_add_66380;
    p32_add_65032 <= p31_add_65032;
    p32_and_66458 <= p32_and_66458_comb;
    p32_add_66479 <= p32_add_66479_comb;
    p32_add_65172 <= p31_add_65172;
  end

  // ===== Pipe stage 33:
  wire [31:0] p33_and_66560_comb;
  wire [31:0] p33_add_66551_comb;
  wire [28:0] p33_add_66556_comb;
  wire [31:0] p33_add_66552_comb;
  wire [31:0] p33_add_66579_comb;
  wire [31:0] p33_add_66553_comb;
  wire [31:0] p33_add_66559_comb;
  wire [31:0] p33_add_66581_comb;
  assign p33_and_66560_comb = p32_add_66479 & p32_add_66380;
  assign p33_add_66551_comb = {p32_add_66454[5:0] ^ p32_add_66454[10:5] ^ p32_add_66454[24:19], p32_add_66454[31:27] ^ p32_add_66454[4:0] ^ p32_add_66454[18:14], p32_add_66454[26:13] ^ p32_add_66454[31:18] ^ p32_add_66454[13:0], p32_add_66454[12:6] ^ p32_add_66454[17:11] ^ p32_add_66454[31:25]} + (p32_add_66454 & p32_add_66355 ^ ~(p32_add_66454 | ~p32_add_66256));
  assign p33_add_66556_comb = p32_add_64891[31:3] + 29'h05c3_6427;
  assign p33_add_66552_comb = p33_add_66551_comb + p32_add_66457;
  assign p33_add_66579_comb = (p33_and_66560_comb ^ p32_add_66479 & p32_add_66281 ^ p32_and_66458) + p32_add_66453;
  assign p33_add_66553_comb = p33_add_66552_comb + p32_add_66281;
  assign p33_add_66559_comb = {p33_add_66556_comb, p32_add_64891[2:0]} + p32_add_66256;
  assign p33_add_66581_comb = p33_add_66579_comb + {p32_add_66479[1:0] ^ p32_add_66479[12:11] ^ p32_add_66479[21:20], p32_add_66479[31:21] ^ p32_add_66479[10:0] ^ p32_add_66479[19:9], p32_add_66479[20:12] ^ p32_add_66479[31:23] ^ p32_add_66479[8:0], p32_add_66479[11:2] ^ p32_add_66479[22:13] ^ p32_add_66479[31:22]};

  // Registers for pipe stage 33:
  reg [31:0] p33_add_63775;
  reg [31:0] p33_add_64102;
  reg [31:0] p33_add_63845;
  reg [31:0] p33_add_64121;
  reg [31:0] p33_add_64138;
  reg [31:0] p33_add_64290;
  reg [31:0] p33_add_64291;
  reg [31:0] p33_add_64441;
  reg [31:0] p33_add_64326;
  reg [31:0] p33_add_64459;
  reg [31:0] p33_add_64477;
  reg [31:0] p33_add_66355;
  reg [31:0] p33_add_64612;
  reg [31:0] p33_add_66454;
  reg [31:0] p33_add_64750;
  reg [31:0] p33_add_66552;
  reg [31:0] p33_add_66553;
  reg [31:0] p33_add_64891;
  reg [31:0] p33_add_66559;
  reg [31:0] p33_add_66380;
  reg [31:0] p33_add_65032;
  reg [31:0] p33_add_66479;
  reg [31:0] p33_add_65172;
  reg [31:0] p33_and_66560;
  reg [31:0] p33_add_66581;
  always_ff @ (posedge clk) begin
    p33_add_63775 <= p32_add_63775;
    p33_add_64102 <= p32_add_64102;
    p33_add_63845 <= p32_add_63845;
    p33_add_64121 <= p32_add_64121;
    p33_add_64138 <= p32_add_64138;
    p33_add_64290 <= p32_add_64290;
    p33_add_64291 <= p32_add_64291;
    p33_add_64441 <= p32_add_64441;
    p33_add_64326 <= p32_add_64326;
    p33_add_64459 <= p32_add_64459;
    p33_add_64477 <= p32_add_64477;
    p33_add_66355 <= p32_add_66355;
    p33_add_64612 <= p32_add_64612;
    p33_add_66454 <= p32_add_66454;
    p33_add_64750 <= p32_add_64750;
    p33_add_66552 <= p33_add_66552_comb;
    p33_add_66553 <= p33_add_66553_comb;
    p33_add_64891 <= p32_add_64891;
    p33_add_66559 <= p33_add_66559_comb;
    p33_add_66380 <= p32_add_66380;
    p33_add_65032 <= p32_add_65032;
    p33_add_66479 <= p32_add_66479;
    p33_add_65172 <= p32_add_65172;
    p33_and_66560 <= p33_and_66560_comb;
    p33_add_66581 <= p33_add_66581_comb;
  end

  // ===== Pipe stage 34:
  wire [31:0] p34_and_66696_comb;
  wire [31:0] p34_add_66653_comb;
  wire [29:0] p34_add_66658_comb;
  wire [31:0] p34_add_66654_comb;
  wire [31:0] p34_add_66693_comb;
  wire [31:0] p34_add_66694_comb;
  wire [31:0] p34_add_66715_comb;
  wire [31:0] p34_add_66750_comb;
  wire [31:0] p34_add_66751_comb;
  wire [31:0] p34_add_66655_comb;
  wire [31:0] p34_add_66661_comb;
  wire [31:0] p34_add_66695_comb;
  wire [31:0] p34_add_66739_comb;
  wire [31:0] p34_add_66752_comb;
  assign p34_and_66696_comb = p33_add_66581 & p33_add_66479;
  assign p34_add_66653_comb = (p33_add_66553 & p33_add_66454 ^ ~(p33_add_66553 | ~p33_add_66355)) + {p33_add_66553[5:0] ^ p33_add_66553[10:5] ^ p33_add_66553[24:19], p33_add_66553[31:27] ^ p33_add_66553[4:0] ^ p33_add_66553[18:14], p33_add_66553[26:13] ^ p33_add_66553[31:18] ^ p33_add_66553[13:0], p33_add_66553[12:6] ^ p33_add_66553[17:11] ^ p33_add_66553[31:25]};
  assign p34_add_66658_comb = p33_add_65032[31:2] + 30'h134b_1b7f;
  assign p34_add_66654_comb = p34_add_66653_comb + p33_add_66559;
  assign p34_add_66693_comb = p33_add_64459 + {p33_add_64102[6:4] ^ p33_add_64102[17:15], p33_add_64102[3:0] ^ p33_add_64102[14:11] ^ p33_add_64102[31:28], p33_add_64102[31:21] ^ p33_add_64102[10:0] ^ p33_add_64102[27:17], p33_add_64102[20:7] ^ p33_add_64102[31:18] ^ p33_add_64102[16:3]};
  assign p34_add_66694_comb = {p33_add_65032[16:7] ^ p33_add_65032[18:9], p33_add_65032[6:0] ^ p33_add_65032[8:2] ^ p33_add_65032[31:25], p33_add_65032[31:30] ^ p33_add_65032[1:0] ^ p33_add_65032[24:23], p33_add_65032[29:17] ^ p33_add_65032[31:19] ^ p33_add_65032[22:10]} + p33_add_63775;
  assign p34_add_66715_comb = (p34_and_66696_comb ^ p33_add_66581 & p33_add_66380 ^ p33_and_66560) + p33_add_66552;
  assign p34_add_66750_comb = p33_add_64477 + {p33_add_63845[6:4] ^ p33_add_63845[17:15], p33_add_63845[3:0] ^ p33_add_63845[14:11] ^ p33_add_63845[31:28], p33_add_63845[31:21] ^ p33_add_63845[10:0] ^ p33_add_63845[27:17], p33_add_63845[20:7] ^ p33_add_63845[31:18] ^ p33_add_63845[16:3]};
  assign p34_add_66751_comb = {p33_add_65172[16:7] ^ p33_add_65172[18:9], p33_add_65172[6:0] ^ p33_add_65172[8:2] ^ p33_add_65172[31:25], p33_add_65172[31:30] ^ p33_add_65172[1:0] ^ p33_add_65172[24:23], p33_add_65172[29:17] ^ p33_add_65172[31:19] ^ p33_add_65172[22:10]} + p33_add_64102;
  assign p34_add_66655_comb = p34_add_66654_comb + p33_add_66380;
  assign p34_add_66661_comb = {p34_add_66658_comb, p33_add_65032[1:0]} + p33_add_66355;
  assign p34_add_66695_comb = p34_add_66693_comb + p34_add_66694_comb;
  assign p34_add_66739_comb = p34_add_66715_comb + {p33_add_66581[1:0] ^ p33_add_66581[12:11] ^ p33_add_66581[21:20], p33_add_66581[31:21] ^ p33_add_66581[10:0] ^ p33_add_66581[19:9], p33_add_66581[20:12] ^ p33_add_66581[31:23] ^ p33_add_66581[8:0], p33_add_66581[11:2] ^ p33_add_66581[22:13] ^ p33_add_66581[31:22]};
  assign p34_add_66752_comb = p34_add_66750_comb + p34_add_66751_comb;

  // Registers for pipe stage 34:
  reg [31:0] p34_add_63845;
  reg [31:0] p34_add_64121;
  reg [31:0] p34_add_64138;
  reg [31:0] p34_add_64290;
  reg [31:0] p34_add_64291;
  reg [31:0] p34_add_64441;
  reg [31:0] p34_add_64326;
  reg [31:0] p34_add_64459;
  reg [31:0] p34_add_64477;
  reg [31:0] p34_add_64612;
  reg [31:0] p34_add_66454;
  reg [31:0] p34_add_64750;
  reg [31:0] p34_add_66553;
  reg [31:0] p34_add_64891;
  reg [31:0] p34_add_66654;
  reg [31:0] p34_add_66655;
  reg [31:0] p34_add_65032;
  reg [31:0] p34_add_66661;
  reg [31:0] p34_add_66479;
  reg [31:0] p34_add_65172;
  reg [31:0] p34_add_66581;
  reg [31:0] p34_add_66695;
  reg [31:0] p34_and_66696;
  reg [31:0] p34_add_66739;
  reg [31:0] p34_add_66752;
  always_ff @ (posedge clk) begin
    p34_add_63845 <= p33_add_63845;
    p34_add_64121 <= p33_add_64121;
    p34_add_64138 <= p33_add_64138;
    p34_add_64290 <= p33_add_64290;
    p34_add_64291 <= p33_add_64291;
    p34_add_64441 <= p33_add_64441;
    p34_add_64326 <= p33_add_64326;
    p34_add_64459 <= p33_add_64459;
    p34_add_64477 <= p33_add_64477;
    p34_add_64612 <= p33_add_64612;
    p34_add_66454 <= p33_add_66454;
    p34_add_64750 <= p33_add_64750;
    p34_add_66553 <= p33_add_66553;
    p34_add_64891 <= p33_add_64891;
    p34_add_66654 <= p34_add_66654_comb;
    p34_add_66655 <= p34_add_66655_comb;
    p34_add_65032 <= p33_add_65032;
    p34_add_66661 <= p34_add_66661_comb;
    p34_add_66479 <= p33_add_66479;
    p34_add_65172 <= p33_add_65172;
    p34_add_66581 <= p33_add_66581;
    p34_add_66695 <= p34_add_66695_comb;
    p34_and_66696 <= p34_and_66696_comb;
    p34_add_66739 <= p34_add_66739_comb;
    p34_add_66752 <= p34_add_66752_comb;
  end

  // ===== Pipe stage 35:
  wire [1:0] p35_bit_slice_66830_comb;
  wire [31:0] p35_add_66884_comb;
  wire [31:0] p35_add_66885_comb;
  wire [31:0] p35_add_66886_comb;
  wire [31:0] p35_and_66831_comb;
  wire [31:0] p35_add_66824_comb;
  wire [31:0] p35_add_66825_comb;
  wire [31:0] p35_add_66828_comb;
  wire [31:0] p35_add_66879_comb;
  wire [31:0] p35_add_66919_comb;
  wire [31:0] p35_add_66920_comb;
  wire [31:0] p35_add_66826_comb;
  wire [31:0] p35_add_66829_comb;
  wire [31:0] p35_add_66883_comb;
  wire [31:0] p35_add_66921_comb;
  wire [31:0] p35_add_66938_comb;
  assign p35_bit_slice_66830_comb = p34_add_66695[1:0];
  assign p35_add_66884_comb = p34_add_64612 + {p34_add_64121[6:4] ^ p34_add_64121[17:15], p34_add_64121[3:0] ^ p34_add_64121[14:11] ^ p34_add_64121[31:28], p34_add_64121[31:21] ^ p34_add_64121[10:0] ^ p34_add_64121[27:17], p34_add_64121[20:7] ^ p34_add_64121[31:18] ^ p34_add_64121[16:3]};
  assign p35_add_66885_comb = {p34_add_66695[16:7] ^ p34_add_66695[18:9], p34_add_66695[6:0] ^ p34_add_66695[8:2] ^ p34_add_66695[31:25], p34_add_66695[31:30] ^ p35_bit_slice_66830_comb ^ p34_add_66695[24:23], p34_add_66695[29:17] ^ p34_add_66695[31:19] ^ p34_add_66695[22:10]} + p34_add_63845;
  assign p35_add_66886_comb = p35_add_66884_comb + p35_add_66885_comb;
  assign p35_and_66831_comb = p34_add_66739 & p34_add_66581;
  assign p35_add_66824_comb = (p34_add_66655 & p34_add_66553 ^ ~(p34_add_66655 | ~p34_add_66454)) + {p34_add_66655[5:0] ^ p34_add_66655[10:5] ^ p34_add_66655[24:19], p34_add_66655[31:27] ^ p34_add_66655[4:0] ^ p34_add_66655[18:14], p34_add_66655[26:13] ^ p34_add_66655[31:18] ^ p34_add_66655[13:0], p34_add_66655[12:6] ^ p34_add_66655[17:11] ^ p34_add_66655[31:25]};
  assign p35_add_66825_comb = p35_add_66824_comb + p34_add_66661;
  assign p35_add_66828_comb = p34_add_65172 + 32'h5338_0d13;
  assign p35_add_66879_comb = (p35_and_66831_comb ^ p34_add_66739 & p34_add_66479 ^ p34_and_66696) + p34_add_66654;
  assign p35_add_66919_comb = p34_add_64750 + {p34_add_64138[6:4] ^ p34_add_64138[17:15], p34_add_64138[3:0] ^ p34_add_64138[14:11] ^ p34_add_64138[31:28], p34_add_64138[31:21] ^ p34_add_64138[10:0] ^ p34_add_64138[27:17], p34_add_64138[20:7] ^ p34_add_64138[31:18] ^ p34_add_64138[16:3]};
  assign p35_add_66920_comb = {p34_add_66752[16:7] ^ p34_add_66752[18:9], p34_add_66752[6:0] ^ p34_add_66752[8:2] ^ p34_add_66752[31:25], p34_add_66752[31:30] ^ p34_add_66752[1:0] ^ p34_add_66752[24:23], p34_add_66752[29:17] ^ p34_add_66752[31:19] ^ p34_add_66752[22:10]} + p34_add_64121;
  assign p35_add_66826_comb = p35_add_66825_comb + p34_add_66479;
  assign p35_add_66829_comb = p34_add_66454 + p35_add_66828_comb;
  assign p35_add_66883_comb = p35_add_66879_comb + {p34_add_66739[1:0] ^ p34_add_66739[12:11] ^ p34_add_66739[21:20], p34_add_66739[31:21] ^ p34_add_66739[10:0] ^ p34_add_66739[19:9], p34_add_66739[20:12] ^ p34_add_66739[31:23] ^ p34_add_66739[8:0], p34_add_66739[11:2] ^ p34_add_66739[22:13] ^ p34_add_66739[31:22]};
  assign p35_add_66921_comb = p35_add_66919_comb + p35_add_66920_comb;
  assign p35_add_66938_comb = {p35_add_66886_comb[16:7] ^ p35_add_66886_comb[18:9], p35_add_66886_comb[6:0] ^ p35_add_66886_comb[8:2] ^ p35_add_66886_comb[31:25], p35_add_66886_comb[31:30] ^ p35_add_66886_comb[1:0] ^ p35_add_66886_comb[24:23], p35_add_66886_comb[29:17] ^ p35_add_66886_comb[31:19] ^ p35_add_66886_comb[22:10]} + p34_add_64138;

  // Registers for pipe stage 35:
  reg [31:0] p35_add_64290;
  reg [31:0] p35_add_64291;
  reg [31:0] p35_add_64441;
  reg [31:0] p35_add_64326;
  reg [31:0] p35_add_64459;
  reg [31:0] p35_add_64477;
  reg [31:0] p35_add_64612;
  reg [31:0] p35_add_64750;
  reg [31:0] p35_add_66553;
  reg [31:0] p35_add_64891;
  reg [31:0] p35_add_66655;
  reg [31:0] p35_add_65032;
  reg [31:0] p35_add_66825;
  reg [31:0] p35_add_66826;
  reg [31:0] p35_add_65172;
  reg [31:0] p35_add_66829;
  reg [31:0] p35_add_66581;
  reg [31:0] p35_add_66695;
  reg [1:0] p35_bit_slice_66830;
  reg [31:0] p35_add_66739;
  reg [31:0] p35_add_66752;
  reg [31:0] p35_and_66831;
  reg [31:0] p35_add_66883;
  reg [31:0] p35_add_66886;
  reg [31:0] p35_add_66921;
  reg [31:0] p35_add_66938;
  always_ff @ (posedge clk) begin
    p35_add_64290 <= p34_add_64290;
    p35_add_64291 <= p34_add_64291;
    p35_add_64441 <= p34_add_64441;
    p35_add_64326 <= p34_add_64326;
    p35_add_64459 <= p34_add_64459;
    p35_add_64477 <= p34_add_64477;
    p35_add_64612 <= p34_add_64612;
    p35_add_64750 <= p34_add_64750;
    p35_add_66553 <= p34_add_66553;
    p35_add_64891 <= p34_add_64891;
    p35_add_66655 <= p34_add_66655;
    p35_add_65032 <= p34_add_65032;
    p35_add_66825 <= p35_add_66825_comb;
    p35_add_66826 <= p35_add_66826_comb;
    p35_add_65172 <= p34_add_65172;
    p35_add_66829 <= p35_add_66829_comb;
    p35_add_66581 <= p34_add_66581;
    p35_add_66695 <= p34_add_66695;
    p35_bit_slice_66830 <= p35_bit_slice_66830_comb;
    p35_add_66739 <= p34_add_66739;
    p35_add_66752 <= p34_add_66752;
    p35_and_66831 <= p35_and_66831_comb;
    p35_add_66883 <= p35_add_66883_comb;
    p35_add_66886 <= p35_add_66886_comb;
    p35_add_66921 <= p35_add_66921_comb;
    p35_add_66938 <= p35_add_66938_comb;
  end

  // ===== Pipe stage 36:
  wire [31:0] p36_add_67058_comb;
  wire [31:0] p36_add_67059_comb;
  wire [31:0] p36_and_67020_comb;
  wire [31:0] p36_add_67012_comb;
  wire [29:0] p36_add_67017_comb;
  wire [31:0] p36_add_67013_comb;
  wire [31:0] p36_add_67039_comb;
  wire [31:0] p36_add_67092_comb;
  wire [31:0] p36_add_67093_comb;
  wire [31:0] p36_add_67014_comb;
  wire [31:0] p36_add_67019_comb;
  wire [31:0] p36_add_67041_comb;
  wire [31:0] p36_add_67094_comb;
  wire [31:0] p36_add_67111_comb;
  assign p36_add_67058_comb = p35_add_64891 + {p35_add_64290[6:4] ^ p35_add_64290[17:15], p35_add_64290[3:0] ^ p35_add_64290[14:11] ^ p35_add_64290[31:28], p35_add_64290[31:21] ^ p35_add_64290[10:0] ^ p35_add_64290[27:17], p35_add_64290[20:7] ^ p35_add_64290[31:18] ^ p35_add_64290[16:3]};
  assign p36_add_67059_comb = p36_add_67058_comb + p35_add_66938;
  assign p36_and_67020_comb = p35_add_66883 & p35_add_66739;
  assign p36_add_67012_comb = {p35_add_66826[5:0] ^ p35_add_66826[10:5] ^ p35_add_66826[24:19], p35_add_66826[31:27] ^ p35_add_66826[4:0] ^ p35_add_66826[18:14], p35_add_66826[26:13] ^ p35_add_66826[31:18] ^ p35_add_66826[13:0], p35_add_66826[12:6] ^ p35_add_66826[17:11] ^ p35_add_66826[31:25]} + (p35_add_66826 & p35_add_66655 ^ ~(p35_add_66826 | ~p35_add_66553));
  assign p36_add_67017_comb = p35_add_66695[31:2] + 30'h1942_9cd5;
  assign p36_add_67013_comb = p36_add_67012_comb + p35_add_66829;
  assign p36_add_67039_comb = (p36_and_67020_comb ^ p35_add_66883 & p35_add_66581 ^ p35_and_66831) + p35_add_66825;
  assign p36_add_67092_comb = p35_add_65032 + {p35_add_64291[6:4] ^ p35_add_64291[17:15], p35_add_64291[3:0] ^ p35_add_64291[14:11] ^ p35_add_64291[31:28], p35_add_64291[31:21] ^ p35_add_64291[10:0] ^ p35_add_64291[27:17], p35_add_64291[20:7] ^ p35_add_64291[31:18] ^ p35_add_64291[16:3]};
  assign p36_add_67093_comb = {p35_add_66921[16:7] ^ p35_add_66921[18:9], p35_add_66921[6:0] ^ p35_add_66921[8:2] ^ p35_add_66921[31:25], p35_add_66921[31:30] ^ p35_add_66921[1:0] ^ p35_add_66921[24:23], p35_add_66921[29:17] ^ p35_add_66921[31:19] ^ p35_add_66921[22:10]} + p35_add_64290;
  assign p36_add_67014_comb = p36_add_67013_comb + p35_add_66581;
  assign p36_add_67019_comb = {p36_add_67017_comb, p35_bit_slice_66830} + p35_add_66553;
  assign p36_add_67041_comb = p36_add_67039_comb + {p35_add_66883[1:0] ^ p35_add_66883[12:11] ^ p35_add_66883[21:20], p35_add_66883[31:21] ^ p35_add_66883[10:0] ^ p35_add_66883[19:9], p35_add_66883[20:12] ^ p35_add_66883[31:23] ^ p35_add_66883[8:0], p35_add_66883[11:2] ^ p35_add_66883[22:13] ^ p35_add_66883[31:22]};
  assign p36_add_67094_comb = p36_add_67092_comb + p36_add_67093_comb;
  assign p36_add_67111_comb = {p36_add_67059_comb[16:7] ^ p36_add_67059_comb[18:9], p36_add_67059_comb[6:0] ^ p36_add_67059_comb[8:2] ^ p36_add_67059_comb[31:25], p36_add_67059_comb[31:30] ^ p36_add_67059_comb[1:0] ^ p36_add_67059_comb[24:23], p36_add_67059_comb[29:17] ^ p36_add_67059_comb[31:19] ^ p36_add_67059_comb[22:10]} + p35_add_64291;

  // Registers for pipe stage 36:
  reg [31:0] p36_add_64441;
  reg [31:0] p36_add_64326;
  reg [31:0] p36_add_64459;
  reg [31:0] p36_add_64477;
  reg [31:0] p36_add_64612;
  reg [31:0] p36_add_64750;
  reg [31:0] p36_add_64891;
  reg [31:0] p36_add_66655;
  reg [31:0] p36_add_65032;
  reg [31:0] p36_add_66826;
  reg [31:0] p36_add_65172;
  reg [31:0] p36_add_67013;
  reg [31:0] p36_add_67014;
  reg [31:0] p36_add_66695;
  reg [31:0] p36_add_67019;
  reg [31:0] p36_add_66739;
  reg [31:0] p36_add_66752;
  reg [31:0] p36_add_66883;
  reg [31:0] p36_add_66886;
  reg [31:0] p36_and_67020;
  reg [31:0] p36_add_67041;
  reg [31:0] p36_add_66921;
  reg [31:0] p36_add_67059;
  reg [31:0] p36_add_67094;
  reg [31:0] p36_add_67111;
  always_ff @ (posedge clk) begin
    p36_add_64441 <= p35_add_64441;
    p36_add_64326 <= p35_add_64326;
    p36_add_64459 <= p35_add_64459;
    p36_add_64477 <= p35_add_64477;
    p36_add_64612 <= p35_add_64612;
    p36_add_64750 <= p35_add_64750;
    p36_add_64891 <= p35_add_64891;
    p36_add_66655 <= p35_add_66655;
    p36_add_65032 <= p35_add_65032;
    p36_add_66826 <= p35_add_66826;
    p36_add_65172 <= p35_add_65172;
    p36_add_67013 <= p36_add_67013_comb;
    p36_add_67014 <= p36_add_67014_comb;
    p36_add_66695 <= p35_add_66695;
    p36_add_67019 <= p36_add_67019_comb;
    p36_add_66739 <= p35_add_66739;
    p36_add_66752 <= p35_add_66752;
    p36_add_66883 <= p35_add_66883;
    p36_add_66886 <= p35_add_66886;
    p36_and_67020 <= p36_and_67020_comb;
    p36_add_67041 <= p36_add_67041_comb;
    p36_add_66921 <= p35_add_66921;
    p36_add_67059 <= p36_add_67059_comb;
    p36_add_67094 <= p36_add_67094_comb;
    p36_add_67111 <= p36_add_67111_comb;
  end

  // ===== Pipe stage 37:
  wire [31:0] p37_add_67227_comb;
  wire [31:0] p37_add_67228_comb;
  wire [31:0] p37_and_67189_comb;
  wire [31:0] p37_add_67183_comb;
  wire [31:0] p37_add_67184_comb;
  wire [31:0] p37_add_67187_comb;
  wire [31:0] p37_add_67208_comb;
  wire [31:0] p37_add_67261_comb;
  wire [31:0] p37_add_67262_comb;
  wire [31:0] p37_add_67185_comb;
  wire [31:0] p37_add_67188_comb;
  wire [31:0] p37_add_67210_comb;
  wire [31:0] p37_add_67263_comb;
  wire [31:0] p37_add_67280_comb;
  assign p37_add_67227_comb = p36_add_65172 + {p36_add_64441[6:4] ^ p36_add_64441[17:15], p36_add_64441[3:0] ^ p36_add_64441[14:11] ^ p36_add_64441[31:28], p36_add_64441[31:21] ^ p36_add_64441[10:0] ^ p36_add_64441[27:17], p36_add_64441[20:7] ^ p36_add_64441[31:18] ^ p36_add_64441[16:3]};
  assign p37_add_67228_comb = p37_add_67227_comb + p36_add_67111;
  assign p37_and_67189_comb = p36_add_67041 & p36_add_66883;
  assign p37_add_67183_comb = (p36_add_67014 & p36_add_66826 ^ ~(p36_add_67014 | ~p36_add_66655)) + {p36_add_67014[5:0] ^ p36_add_67014[10:5] ^ p36_add_67014[24:19], p36_add_67014[31:27] ^ p36_add_67014[4:0] ^ p36_add_67014[18:14], p36_add_67014[26:13] ^ p36_add_67014[31:18] ^ p36_add_67014[13:0], p36_add_67014[12:6] ^ p36_add_67014[17:11] ^ p36_add_67014[31:25]};
  assign p37_add_67184_comb = p37_add_67183_comb + p36_add_67019;
  assign p37_add_67187_comb = p36_add_66752 + 32'h766a_0abb;
  assign p37_add_67208_comb = (p37_and_67189_comb ^ p36_add_67041 & p36_add_66739 ^ p36_and_67020) + p36_add_67013;
  assign p37_add_67261_comb = p36_add_66695 + {p36_add_64326[6:4] ^ p36_add_64326[17:15], p36_add_64326[3:0] ^ p36_add_64326[14:11] ^ p36_add_64326[31:28], p36_add_64326[31:21] ^ p36_add_64326[10:0] ^ p36_add_64326[27:17], p36_add_64326[20:7] ^ p36_add_64326[31:18] ^ p36_add_64326[16:3]};
  assign p37_add_67262_comb = {p36_add_67094[16:7] ^ p36_add_67094[18:9], p36_add_67094[6:0] ^ p36_add_67094[8:2] ^ p36_add_67094[31:25], p36_add_67094[31:30] ^ p36_add_67094[1:0] ^ p36_add_67094[24:23], p36_add_67094[29:17] ^ p36_add_67094[31:19] ^ p36_add_67094[22:10]} + p36_add_64441;
  assign p37_add_67185_comb = p37_add_67184_comb + p36_add_66739;
  assign p37_add_67188_comb = p36_add_66655 + p37_add_67187_comb;
  assign p37_add_67210_comb = p37_add_67208_comb + {p36_add_67041[1:0] ^ p36_add_67041[12:11] ^ p36_add_67041[21:20], p36_add_67041[31:21] ^ p36_add_67041[10:0] ^ p36_add_67041[19:9], p36_add_67041[20:12] ^ p36_add_67041[31:23] ^ p36_add_67041[8:0], p36_add_67041[11:2] ^ p36_add_67041[22:13] ^ p36_add_67041[31:22]};
  assign p37_add_67263_comb = p37_add_67261_comb + p37_add_67262_comb;
  assign p37_add_67280_comb = {p37_add_67228_comb[16:7] ^ p37_add_67228_comb[18:9], p37_add_67228_comb[6:0] ^ p37_add_67228_comb[8:2] ^ p37_add_67228_comb[31:25], p37_add_67228_comb[31:30] ^ p37_add_67228_comb[1:0] ^ p37_add_67228_comb[24:23], p37_add_67228_comb[29:17] ^ p37_add_67228_comb[31:19] ^ p37_add_67228_comb[22:10]} + p36_add_64326;

  // Registers for pipe stage 37:
  reg [31:0] p37_add_64459;
  reg [31:0] p37_add_64477;
  reg [31:0] p37_add_64612;
  reg [31:0] p37_add_64750;
  reg [31:0] p37_add_64891;
  reg [31:0] p37_add_65032;
  reg [31:0] p37_add_66826;
  reg [31:0] p37_add_65172;
  reg [31:0] p37_add_67014;
  reg [31:0] p37_add_66695;
  reg [31:0] p37_add_67184;
  reg [31:0] p37_add_67185;
  reg [31:0] p37_add_66752;
  reg [31:0] p37_add_67188;
  reg [31:0] p37_add_66883;
  reg [31:0] p37_add_66886;
  reg [31:0] p37_add_67041;
  reg [31:0] p37_add_66921;
  reg [31:0] p37_and_67189;
  reg [31:0] p37_add_67210;
  reg [31:0] p37_add_67059;
  reg [31:0] p37_add_67094;
  reg [31:0] p37_add_67228;
  reg [31:0] p37_add_67263;
  reg [31:0] p37_add_67280;
  always_ff @ (posedge clk) begin
    p37_add_64459 <= p36_add_64459;
    p37_add_64477 <= p36_add_64477;
    p37_add_64612 <= p36_add_64612;
    p37_add_64750 <= p36_add_64750;
    p37_add_64891 <= p36_add_64891;
    p37_add_65032 <= p36_add_65032;
    p37_add_66826 <= p36_add_66826;
    p37_add_65172 <= p36_add_65172;
    p37_add_67014 <= p36_add_67014;
    p37_add_66695 <= p36_add_66695;
    p37_add_67184 <= p37_add_67184_comb;
    p37_add_67185 <= p37_add_67185_comb;
    p37_add_66752 <= p36_add_66752;
    p37_add_67188 <= p37_add_67188_comb;
    p37_add_66883 <= p36_add_66883;
    p37_add_66886 <= p36_add_66886;
    p37_add_67041 <= p36_add_67041;
    p37_add_66921 <= p36_add_66921;
    p37_and_67189 <= p37_and_67189_comb;
    p37_add_67210 <= p37_add_67210_comb;
    p37_add_67059 <= p36_add_67059;
    p37_add_67094 <= p36_add_67094;
    p37_add_67228 <= p37_add_67228_comb;
    p37_add_67263 <= p37_add_67263_comb;
    p37_add_67280 <= p37_add_67280_comb;
  end

  // ===== Pipe stage 38:
  wire [31:0] p38_add_67399_comb;
  wire [31:0] p38_add_67400_comb;
  wire [31:0] p38_and_67361_comb;
  wire [31:0] p38_add_67352_comb;
  wire [30:0] p38_add_67357_comb;
  wire [31:0] p38_add_67353_comb;
  wire [31:0] p38_add_67380_comb;
  wire [31:0] p38_add_67433_comb;
  wire [31:0] p38_add_67434_comb;
  wire [31:0] p38_add_67354_comb;
  wire [31:0] p38_add_67360_comb;
  wire [31:0] p38_add_67382_comb;
  wire [31:0] p38_add_67435_comb;
  wire [31:0] p38_add_67452_comb;
  assign p38_add_67399_comb = p37_add_66752 + {p37_add_64459[6:4] ^ p37_add_64459[17:15], p37_add_64459[3:0] ^ p37_add_64459[14:11] ^ p37_add_64459[31:28], p37_add_64459[31:21] ^ p37_add_64459[10:0] ^ p37_add_64459[27:17], p37_add_64459[20:7] ^ p37_add_64459[31:18] ^ p37_add_64459[16:3]};
  assign p38_add_67400_comb = p38_add_67399_comb + p37_add_67280;
  assign p38_and_67361_comb = p37_add_67210 & p37_add_67041;
  assign p38_add_67352_comb = {p37_add_67185[5:0] ^ p37_add_67185[10:5] ^ p37_add_67185[24:19], p37_add_67185[31:27] ^ p37_add_67185[4:0] ^ p37_add_67185[18:14], p37_add_67185[26:13] ^ p37_add_67185[31:18] ^ p37_add_67185[13:0], p37_add_67185[12:6] ^ p37_add_67185[17:11] ^ p37_add_67185[31:25]} + (p37_add_67185 & p37_add_67014 ^ ~(p37_add_67185 | ~p37_add_66826));
  assign p38_add_67357_comb = p37_add_66886[31:1] + 31'h40e1_6497;
  assign p38_add_67353_comb = p38_add_67352_comb + p37_add_67188;
  assign p38_add_67380_comb = (p38_and_67361_comb ^ p37_add_67210 & p37_add_66883 ^ p37_and_67189) + p37_add_67184;
  assign p38_add_67433_comb = p37_add_66886 + {p37_add_64477[6:4] ^ p37_add_64477[17:15], p37_add_64477[3:0] ^ p37_add_64477[14:11] ^ p37_add_64477[31:28], p37_add_64477[31:21] ^ p37_add_64477[10:0] ^ p37_add_64477[27:17], p37_add_64477[20:7] ^ p37_add_64477[31:18] ^ p37_add_64477[16:3]};
  assign p38_add_67434_comb = {p37_add_67263[16:7] ^ p37_add_67263[18:9], p37_add_67263[6:0] ^ p37_add_67263[8:2] ^ p37_add_67263[31:25], p37_add_67263[31:30] ^ p37_add_67263[1:0] ^ p37_add_67263[24:23], p37_add_67263[29:17] ^ p37_add_67263[31:19] ^ p37_add_67263[22:10]} + p37_add_64459;
  assign p38_add_67354_comb = p38_add_67353_comb + p37_add_66883;
  assign p38_add_67360_comb = {p38_add_67357_comb, p37_add_66886[0]} + p37_add_66826;
  assign p38_add_67382_comb = p38_add_67380_comb + {p37_add_67210[1:0] ^ p37_add_67210[12:11] ^ p37_add_67210[21:20], p37_add_67210[31:21] ^ p37_add_67210[10:0] ^ p37_add_67210[19:9], p37_add_67210[20:12] ^ p37_add_67210[31:23] ^ p37_add_67210[8:0], p37_add_67210[11:2] ^ p37_add_67210[22:13] ^ p37_add_67210[31:22]};
  assign p38_add_67435_comb = p38_add_67433_comb + p38_add_67434_comb;
  assign p38_add_67452_comb = {p38_add_67400_comb[16:7] ^ p38_add_67400_comb[18:9], p38_add_67400_comb[6:0] ^ p38_add_67400_comb[8:2] ^ p38_add_67400_comb[31:25], p38_add_67400_comb[31:30] ^ p38_add_67400_comb[1:0] ^ p38_add_67400_comb[24:23], p38_add_67400_comb[29:17] ^ p38_add_67400_comb[31:19] ^ p38_add_67400_comb[22:10]} + p37_add_64477;

  // Registers for pipe stage 38:
  reg [31:0] p38_add_64612;
  reg [31:0] p38_add_64750;
  reg [31:0] p38_add_64891;
  reg [31:0] p38_add_65032;
  reg [31:0] p38_add_65172;
  reg [31:0] p38_add_67014;
  reg [31:0] p38_add_66695;
  reg [31:0] p38_add_67185;
  reg [31:0] p38_add_66752;
  reg [31:0] p38_add_67353;
  reg [31:0] p38_add_67354;
  reg [31:0] p38_add_66886;
  reg [31:0] p38_add_67360;
  reg [31:0] p38_add_67041;
  reg [31:0] p38_add_66921;
  reg [31:0] p38_add_67210;
  reg [31:0] p38_add_67059;
  reg [31:0] p38_and_67361;
  reg [31:0] p38_add_67382;
  reg [31:0] p38_add_67094;
  reg [31:0] p38_add_67228;
  reg [31:0] p38_add_67263;
  reg [31:0] p38_add_67400;
  reg [31:0] p38_add_67435;
  reg [31:0] p38_add_67452;
  always_ff @ (posedge clk) begin
    p38_add_64612 <= p37_add_64612;
    p38_add_64750 <= p37_add_64750;
    p38_add_64891 <= p37_add_64891;
    p38_add_65032 <= p37_add_65032;
    p38_add_65172 <= p37_add_65172;
    p38_add_67014 <= p37_add_67014;
    p38_add_66695 <= p37_add_66695;
    p38_add_67185 <= p37_add_67185;
    p38_add_66752 <= p37_add_66752;
    p38_add_67353 <= p38_add_67353_comb;
    p38_add_67354 <= p38_add_67354_comb;
    p38_add_66886 <= p37_add_66886;
    p38_add_67360 <= p38_add_67360_comb;
    p38_add_67041 <= p37_add_67041;
    p38_add_66921 <= p37_add_66921;
    p38_add_67210 <= p37_add_67210;
    p38_add_67059 <= p37_add_67059;
    p38_and_67361 <= p38_and_67361_comb;
    p38_add_67382 <= p38_add_67382_comb;
    p38_add_67094 <= p37_add_67094;
    p38_add_67228 <= p37_add_67228;
    p38_add_67263 <= p37_add_67263;
    p38_add_67400 <= p38_add_67400_comb;
    p38_add_67435 <= p38_add_67435_comb;
    p38_add_67452 <= p38_add_67452_comb;
  end

  // ===== Pipe stage 39:
  wire [31:0] p39_add_67569_comb;
  wire [1:0] p39_bit_slice_67552_comb;
  wire [31:0] p39_add_67570_comb;
  wire [31:0] p39_and_67530_comb;
  wire [31:0] p39_add_67524_comb;
  wire [31:0] p39_add_67525_comb;
  wire [31:0] p39_add_67528_comb;
  wire [31:0] p39_add_67549_comb;
  wire [31:0] p39_add_67602_comb;
  wire [31:0] p39_add_67603_comb;
  wire [31:0] p39_add_67526_comb;
  wire [31:0] p39_add_67529_comb;
  wire [31:0] p39_add_67551_comb;
  wire [31:0] p39_add_67604_comb;
  wire [31:0] p39_add_67621_comb;
  assign p39_add_67569_comb = p38_add_66921 + {p38_add_64612[6:4] ^ p38_add_64612[17:15], p38_add_64612[3:0] ^ p38_add_64612[14:11] ^ p38_add_64612[31:28], p38_add_64612[31:21] ^ p38_add_64612[10:0] ^ p38_add_64612[27:17], p38_add_64612[20:7] ^ p38_add_64612[31:18] ^ p38_add_64612[16:3]};
  assign p39_bit_slice_67552_comb = p38_add_67435[1:0];
  assign p39_add_67570_comb = p39_add_67569_comb + p38_add_67452;
  assign p39_and_67530_comb = p38_add_67382 & p38_add_67210;
  assign p39_add_67524_comb = (p38_add_67354 & p38_add_67185 ^ ~(p38_add_67354 | ~p38_add_67014)) + {p38_add_67354[5:0] ^ p38_add_67354[10:5] ^ p38_add_67354[24:19], p38_add_67354[31:27] ^ p38_add_67354[4:0] ^ p38_add_67354[18:14], p38_add_67354[26:13] ^ p38_add_67354[31:18] ^ p38_add_67354[13:0], p38_add_67354[12:6] ^ p38_add_67354[17:11] ^ p38_add_67354[31:25]};
  assign p39_add_67525_comb = p39_add_67524_comb + p38_add_67360;
  assign p39_add_67528_comb = p38_add_66921 + 32'h9272_2c85;
  assign p39_add_67549_comb = (p39_and_67530_comb ^ p38_add_67382 & p38_add_67041 ^ p38_and_67361) + p38_add_67353;
  assign p39_add_67602_comb = p38_add_67059 + {p38_add_64750[6:4] ^ p38_add_64750[17:15], p38_add_64750[3:0] ^ p38_add_64750[14:11] ^ p38_add_64750[31:28], p38_add_64750[31:21] ^ p38_add_64750[10:0] ^ p38_add_64750[27:17], p38_add_64750[20:7] ^ p38_add_64750[31:18] ^ p38_add_64750[16:3]};
  assign p39_add_67603_comb = {p38_add_67435[16:7] ^ p38_add_67435[18:9], p38_add_67435[6:0] ^ p38_add_67435[8:2] ^ p38_add_67435[31:25], p38_add_67435[31:30] ^ p39_bit_slice_67552_comb ^ p38_add_67435[24:23], p38_add_67435[29:17] ^ p38_add_67435[31:19] ^ p38_add_67435[22:10]} + p38_add_64612;
  assign p39_add_67526_comb = p39_add_67525_comb + p38_add_67041;
  assign p39_add_67529_comb = p38_add_67014 + p39_add_67528_comb;
  assign p39_add_67551_comb = p39_add_67549_comb + {p38_add_67382[1:0] ^ p38_add_67382[12:11] ^ p38_add_67382[21:20], p38_add_67382[31:21] ^ p38_add_67382[10:0] ^ p38_add_67382[19:9], p38_add_67382[20:12] ^ p38_add_67382[31:23] ^ p38_add_67382[8:0], p38_add_67382[11:2] ^ p38_add_67382[22:13] ^ p38_add_67382[31:22]};
  assign p39_add_67604_comb = p39_add_67602_comb + p39_add_67603_comb;
  assign p39_add_67621_comb = {p39_add_67570_comb[16:7] ^ p39_add_67570_comb[18:9], p39_add_67570_comb[6:0] ^ p39_add_67570_comb[8:2] ^ p39_add_67570_comb[31:25], p39_add_67570_comb[31:30] ^ p39_add_67570_comb[1:0] ^ p39_add_67570_comb[24:23], p39_add_67570_comb[29:17] ^ p39_add_67570_comb[31:19] ^ p39_add_67570_comb[22:10]} + p38_add_64750;

  // Registers for pipe stage 39:
  reg [31:0] p39_add_64891;
  reg [31:0] p39_add_65032;
  reg [31:0] p39_add_65172;
  reg [31:0] p39_add_66695;
  reg [31:0] p39_add_67185;
  reg [31:0] p39_add_66752;
  reg [31:0] p39_add_67354;
  reg [31:0] p39_add_66886;
  reg [31:0] p39_add_67525;
  reg [31:0] p39_add_67526;
  reg [31:0] p39_add_66921;
  reg [31:0] p39_add_67529;
  reg [31:0] p39_add_67210;
  reg [31:0] p39_add_67059;
  reg [31:0] p39_add_67382;
  reg [31:0] p39_add_67094;
  reg [31:0] p39_and_67530;
  reg [31:0] p39_add_67551;
  reg [31:0] p39_add_67228;
  reg [31:0] p39_add_67263;
  reg [31:0] p39_add_67400;
  reg [31:0] p39_add_67435;
  reg [1:0] p39_bit_slice_67552;
  reg [31:0] p39_add_67570;
  reg [31:0] p39_add_67604;
  reg [31:0] p39_add_67621;
  always_ff @ (posedge clk) begin
    p39_add_64891 <= p38_add_64891;
    p39_add_65032 <= p38_add_65032;
    p39_add_65172 <= p38_add_65172;
    p39_add_66695 <= p38_add_66695;
    p39_add_67185 <= p38_add_67185;
    p39_add_66752 <= p38_add_66752;
    p39_add_67354 <= p38_add_67354;
    p39_add_66886 <= p38_add_66886;
    p39_add_67525 <= p39_add_67525_comb;
    p39_add_67526 <= p39_add_67526_comb;
    p39_add_66921 <= p38_add_66921;
    p39_add_67529 <= p39_add_67529_comb;
    p39_add_67210 <= p38_add_67210;
    p39_add_67059 <= p38_add_67059;
    p39_add_67382 <= p38_add_67382;
    p39_add_67094 <= p38_add_67094;
    p39_and_67530 <= p39_and_67530_comb;
    p39_add_67551 <= p39_add_67551_comb;
    p39_add_67228 <= p38_add_67228;
    p39_add_67263 <= p38_add_67263;
    p39_add_67400 <= p38_add_67400;
    p39_add_67435 <= p38_add_67435;
    p39_bit_slice_67552 <= p39_bit_slice_67552_comb;
    p39_add_67570 <= p39_add_67570_comb;
    p39_add_67604 <= p39_add_67604_comb;
    p39_add_67621 <= p39_add_67621_comb;
  end

  // ===== Pipe stage 40:
  wire [31:0] p40_add_67739_comb;
  wire [31:0] p40_add_67740_comb;
  wire [31:0] p40_and_67701_comb;
  wire [31:0] p40_add_67695_comb;
  wire [31:0] p40_add_67696_comb;
  wire [31:0] p40_add_67699_comb;
  wire [31:0] p40_add_67720_comb;
  wire [31:0] p40_add_67773_comb;
  wire [31:0] p40_add_67774_comb;
  wire [31:0] p40_add_67697_comb;
  wire [31:0] p40_add_67700_comb;
  wire [31:0] p40_add_67722_comb;
  wire [31:0] p40_add_67775_comb;
  wire [31:0] p40_add_67792_comb;
  assign p40_add_67739_comb = p39_add_67094 + {p39_add_64891[6:4] ^ p39_add_64891[17:15], p39_add_64891[3:0] ^ p39_add_64891[14:11] ^ p39_add_64891[31:28], p39_add_64891[31:21] ^ p39_add_64891[10:0] ^ p39_add_64891[27:17], p39_add_64891[20:7] ^ p39_add_64891[31:18] ^ p39_add_64891[16:3]};
  assign p40_add_67740_comb = p40_add_67739_comb + p39_add_67621;
  assign p40_and_67701_comb = p39_add_67551 & p39_add_67382;
  assign p40_add_67695_comb = {p39_add_67526[5:0] ^ p39_add_67526[10:5] ^ p39_add_67526[24:19], p39_add_67526[31:27] ^ p39_add_67526[4:0] ^ p39_add_67526[18:14], p39_add_67526[26:13] ^ p39_add_67526[31:18] ^ p39_add_67526[13:0], p39_add_67526[12:6] ^ p39_add_67526[17:11] ^ p39_add_67526[31:25]} + (p39_add_67526 & p39_add_67354 ^ ~(p39_add_67526 | ~p39_add_67185));
  assign p40_add_67696_comb = p40_add_67695_comb + p39_add_67529;
  assign p40_add_67699_comb = p39_add_67059 + 32'ha2bf_e8a1;
  assign p40_add_67720_comb = (p40_and_67701_comb ^ p39_add_67551 & p39_add_67210 ^ p39_and_67530) + p39_add_67525;
  assign p40_add_67773_comb = p39_add_67228 + {p39_add_65032[6:4] ^ p39_add_65032[17:15], p39_add_65032[3:0] ^ p39_add_65032[14:11] ^ p39_add_65032[31:28], p39_add_65032[31:21] ^ p39_add_65032[10:0] ^ p39_add_65032[27:17], p39_add_65032[20:7] ^ p39_add_65032[31:18] ^ p39_add_65032[16:3]};
  assign p40_add_67774_comb = {p39_add_67604[16:7] ^ p39_add_67604[18:9], p39_add_67604[6:0] ^ p39_add_67604[8:2] ^ p39_add_67604[31:25], p39_add_67604[31:30] ^ p39_add_67604[1:0] ^ p39_add_67604[24:23], p39_add_67604[29:17] ^ p39_add_67604[31:19] ^ p39_add_67604[22:10]} + p39_add_64891;
  assign p40_add_67697_comb = p40_add_67696_comb + p39_add_67210;
  assign p40_add_67700_comb = p39_add_67185 + p40_add_67699_comb;
  assign p40_add_67722_comb = p40_add_67720_comb + {p39_add_67551[1:0] ^ p39_add_67551[12:11] ^ p39_add_67551[21:20], p39_add_67551[31:21] ^ p39_add_67551[10:0] ^ p39_add_67551[19:9], p39_add_67551[20:12] ^ p39_add_67551[31:23] ^ p39_add_67551[8:0], p39_add_67551[11:2] ^ p39_add_67551[22:13] ^ p39_add_67551[31:22]};
  assign p40_add_67775_comb = p40_add_67773_comb + p40_add_67774_comb;
  assign p40_add_67792_comb = {p40_add_67740_comb[16:7] ^ p40_add_67740_comb[18:9], p40_add_67740_comb[6:0] ^ p40_add_67740_comb[8:2] ^ p40_add_67740_comb[31:25], p40_add_67740_comb[31:30] ^ p40_add_67740_comb[1:0] ^ p40_add_67740_comb[24:23], p40_add_67740_comb[29:17] ^ p40_add_67740_comb[31:19] ^ p40_add_67740_comb[22:10]} + p39_add_65032;

  // Registers for pipe stage 40:
  reg [31:0] p40_add_65172;
  reg [31:0] p40_add_66695;
  reg [31:0] p40_add_66752;
  reg [31:0] p40_add_67354;
  reg [31:0] p40_add_66886;
  reg [31:0] p40_add_67526;
  reg [31:0] p40_add_66921;
  reg [31:0] p40_add_67696;
  reg [31:0] p40_add_67697;
  reg [31:0] p40_add_67059;
  reg [31:0] p40_add_67700;
  reg [31:0] p40_add_67382;
  reg [31:0] p40_add_67094;
  reg [31:0] p40_add_67551;
  reg [31:0] p40_add_67228;
  reg [31:0] p40_and_67701;
  reg [31:0] p40_add_67722;
  reg [31:0] p40_add_67263;
  reg [31:0] p40_add_67400;
  reg [31:0] p40_add_67435;
  reg [1:0] p40_bit_slice_67552;
  reg [31:0] p40_add_67570;
  reg [31:0] p40_add_67604;
  reg [31:0] p40_add_67740;
  reg [31:0] p40_add_67775;
  reg [31:0] p40_add_67792;
  always_ff @ (posedge clk) begin
    p40_add_65172 <= p39_add_65172;
    p40_add_66695 <= p39_add_66695;
    p40_add_66752 <= p39_add_66752;
    p40_add_67354 <= p39_add_67354;
    p40_add_66886 <= p39_add_66886;
    p40_add_67526 <= p39_add_67526;
    p40_add_66921 <= p39_add_66921;
    p40_add_67696 <= p40_add_67696_comb;
    p40_add_67697 <= p40_add_67697_comb;
    p40_add_67059 <= p39_add_67059;
    p40_add_67700 <= p40_add_67700_comb;
    p40_add_67382 <= p39_add_67382;
    p40_add_67094 <= p39_add_67094;
    p40_add_67551 <= p39_add_67551;
    p40_add_67228 <= p39_add_67228;
    p40_and_67701 <= p40_and_67701_comb;
    p40_add_67722 <= p40_add_67722_comb;
    p40_add_67263 <= p39_add_67263;
    p40_add_67400 <= p39_add_67400;
    p40_add_67435 <= p39_add_67435;
    p40_bit_slice_67552 <= p39_bit_slice_67552;
    p40_add_67570 <= p39_add_67570;
    p40_add_67604 <= p39_add_67604;
    p40_add_67740 <= p40_add_67740_comb;
    p40_add_67775 <= p40_add_67775_comb;
    p40_add_67792 <= p40_add_67792_comb;
  end

  // ===== Pipe stage 41:
  wire [31:0] p41_and_67872_comb;
  wire [31:0] p41_add_67866_comb;
  wire [31:0] p41_add_67867_comb;
  wire [31:0] p41_add_67870_comb;
  wire [31:0] p41_add_67891_comb;
  wire [31:0] p41_add_67910_comb;
  wire [31:0] p41_add_67944_comb;
  wire [31:0] p41_add_67945_comb;
  wire [31:0] p41_add_67868_comb;
  wire [31:0] p41_add_67871_comb;
  wire [31:0] p41_add_67893_comb;
  wire [31:0] p41_add_67911_comb;
  wire [31:0] p41_add_67946_comb;
  assign p41_and_67872_comb = p40_add_67722 & p40_add_67551;
  assign p41_add_67866_comb = {p40_add_67697[5:0] ^ p40_add_67697[10:5] ^ p40_add_67697[24:19], p40_add_67697[31:27] ^ p40_add_67697[4:0] ^ p40_add_67697[18:14], p40_add_67697[26:13] ^ p40_add_67697[31:18] ^ p40_add_67697[13:0], p40_add_67697[12:6] ^ p40_add_67697[17:11] ^ p40_add_67697[31:25]} + (p40_add_67697 & p40_add_67526 ^ ~(p40_add_67697 | ~p40_add_67354));
  assign p41_add_67867_comb = p41_add_67866_comb + p40_add_67700;
  assign p41_add_67870_comb = p40_add_67094 + 32'ha81a_664b;
  assign p41_add_67891_comb = (p41_and_67872_comb ^ p40_add_67722 & p40_add_67382 ^ p40_and_67701) + p40_add_67696;
  assign p41_add_67910_comb = p40_add_67263 + {p40_add_65172[6:4] ^ p40_add_65172[17:15], p40_add_65172[3:0] ^ p40_add_65172[14:11] ^ p40_add_65172[31:28], p40_add_65172[31:21] ^ p40_add_65172[10:0] ^ p40_add_65172[27:17], p40_add_65172[20:7] ^ p40_add_65172[31:18] ^ p40_add_65172[16:3]};
  assign p41_add_67944_comb = p40_add_67400 + {p40_add_66695[6:4] ^ p40_add_66695[17:15], p40_add_66695[3:0] ^ p40_add_66695[14:11] ^ p40_add_66695[31:28], p40_add_66695[31:21] ^ p40_add_66695[10:0] ^ p40_add_66695[27:17], p40_add_66695[20:7] ^ p40_add_66695[31:18] ^ p40_add_66695[16:3]};
  assign p41_add_67945_comb = {p40_add_67775[16:7] ^ p40_add_67775[18:9], p40_add_67775[6:0] ^ p40_add_67775[8:2] ^ p40_add_67775[31:25], p40_add_67775[31:30] ^ p40_add_67775[1:0] ^ p40_add_67775[24:23], p40_add_67775[29:17] ^ p40_add_67775[31:19] ^ p40_add_67775[22:10]} + p40_add_65172;
  assign p41_add_67868_comb = p41_add_67867_comb + p40_add_67382;
  assign p41_add_67871_comb = p40_add_67354 + p41_add_67870_comb;
  assign p41_add_67893_comb = p41_add_67891_comb + {p40_add_67722[1:0] ^ p40_add_67722[12:11] ^ p40_add_67722[21:20], p40_add_67722[31:21] ^ p40_add_67722[10:0] ^ p40_add_67722[19:9], p40_add_67722[20:12] ^ p40_add_67722[31:23] ^ p40_add_67722[8:0], p40_add_67722[11:2] ^ p40_add_67722[22:13] ^ p40_add_67722[31:22]};
  assign p41_add_67911_comb = p41_add_67910_comb + p40_add_67792;
  assign p41_add_67946_comb = p41_add_67944_comb + p41_add_67945_comb;

  // Registers for pipe stage 41:
  reg [31:0] p41_add_66695;
  reg [31:0] p41_add_66752;
  reg [31:0] p41_add_66886;
  reg [31:0] p41_add_67526;
  reg [31:0] p41_add_66921;
  reg [31:0] p41_add_67697;
  reg [31:0] p41_add_67059;
  reg [31:0] p41_add_67867;
  reg [31:0] p41_add_67868;
  reg [31:0] p41_add_67094;
  reg [31:0] p41_add_67871;
  reg [31:0] p41_add_67551;
  reg [31:0] p41_add_67228;
  reg [31:0] p41_add_67722;
  reg [31:0] p41_add_67263;
  reg [31:0] p41_and_67872;
  reg [31:0] p41_add_67893;
  reg [31:0] p41_add_67400;
  reg [31:0] p41_add_67435;
  reg [1:0] p41_bit_slice_67552;
  reg [31:0] p41_add_67570;
  reg [31:0] p41_add_67604;
  reg [31:0] p41_add_67740;
  reg [31:0] p41_add_67775;
  reg [31:0] p41_add_67911;
  reg [31:0] p41_add_67946;
  always_ff @ (posedge clk) begin
    p41_add_66695 <= p40_add_66695;
    p41_add_66752 <= p40_add_66752;
    p41_add_66886 <= p40_add_66886;
    p41_add_67526 <= p40_add_67526;
    p41_add_66921 <= p40_add_66921;
    p41_add_67697 <= p40_add_67697;
    p41_add_67059 <= p40_add_67059;
    p41_add_67867 <= p41_add_67867_comb;
    p41_add_67868 <= p41_add_67868_comb;
    p41_add_67094 <= p40_add_67094;
    p41_add_67871 <= p41_add_67871_comb;
    p41_add_67551 <= p40_add_67551;
    p41_add_67228 <= p40_add_67228;
    p41_add_67722 <= p40_add_67722;
    p41_add_67263 <= p40_add_67263;
    p41_and_67872 <= p41_and_67872_comb;
    p41_add_67893 <= p41_add_67893_comb;
    p41_add_67400 <= p40_add_67400;
    p41_add_67435 <= p40_add_67435;
    p41_bit_slice_67552 <= p40_bit_slice_67552;
    p41_add_67570 <= p40_add_67570;
    p41_add_67604 <= p40_add_67604;
    p41_add_67740 <= p40_add_67740;
    p41_add_67775 <= p40_add_67775;
    p41_add_67911 <= p41_add_67911_comb;
    p41_add_67946 <= p41_add_67946_comb;
  end

  // ===== Pipe stage 42:
  wire [1:0] p42_bit_slice_68051_comb;
  wire [31:0] p42_add_68083_comb;
  wire [31:0] p42_add_68084_comb;
  wire [31:0] p42_add_68085_comb;
  wire [31:0] p42_and_68029_comb;
  wire [31:0] p42_add_68020_comb;
  wire [27:0] p42_add_68025_comb;
  wire [31:0] p42_add_68021_comb;
  wire [31:0] p42_add_68048_comb;
  wire [31:0] p42_add_68118_comb;
  wire [31:0] p42_add_68119_comb;
  wire [31:0] p42_add_68022_comb;
  wire [31:0] p42_add_68028_comb;
  wire [31:0] p42_add_68050_comb;
  wire [31:0] p42_add_68120_comb;
  wire [31:0] p42_add_68137_comb;
  wire [3:0] p42_xor_68140_comb;
  assign p42_bit_slice_68051_comb = p41_add_67911[1:0];
  assign p42_add_68083_comb = p41_add_67435 + {p41_add_66752[6:4] ^ p41_add_66752[17:15], p41_add_66752[3:0] ^ p41_add_66752[14:11] ^ p41_add_66752[31:28], p41_add_66752[31:21] ^ p41_add_66752[10:0] ^ p41_add_66752[27:17], p41_add_66752[20:7] ^ p41_add_66752[31:18] ^ p41_add_66752[16:3]};
  assign p42_add_68084_comb = {p41_add_67911[16:7] ^ p41_add_67911[18:9], p41_add_67911[6:0] ^ p41_add_67911[8:2] ^ p41_add_67911[31:25], p41_add_67911[31:30] ^ p42_bit_slice_68051_comb ^ p41_add_67911[24:23], p41_add_67911[29:17] ^ p41_add_67911[31:19] ^ p41_add_67911[22:10]} + p41_add_66695;
  assign p42_add_68085_comb = p42_add_68083_comb + p42_add_68084_comb;
  assign p42_and_68029_comb = p41_add_67893 & p41_add_67722;
  assign p42_add_68020_comb = {p41_add_67868[5:0] ^ p41_add_67868[10:5] ^ p41_add_67868[24:19], p41_add_67868[31:27] ^ p41_add_67868[4:0] ^ p41_add_67868[18:14], p41_add_67868[26:13] ^ p41_add_67868[31:18] ^ p41_add_67868[13:0], p41_add_67868[12:6] ^ p41_add_67868[17:11] ^ p41_add_67868[31:25]} + (p41_add_67868 & p41_add_67697 ^ ~(p41_add_67868 | ~p41_add_67526));
  assign p42_add_68025_comb = p41_add_67228[31:4] + 28'hc24_b8b7;
  assign p42_add_68021_comb = p42_add_68020_comb + p41_add_67871;
  assign p42_add_68048_comb = (p42_and_68029_comb ^ p41_add_67893 & p41_add_67551 ^ p41_and_67872) + p41_add_67867;
  assign p42_add_68118_comb = p41_add_67570 + {p41_add_66886[6:4] ^ p41_add_66886[17:15], p41_add_66886[3:0] ^ p41_add_66886[14:11] ^ p41_add_66886[31:28], p41_add_66886[31:21] ^ p41_add_66886[10:0] ^ p41_add_66886[27:17], p41_add_66886[20:7] ^ p41_add_66886[31:18] ^ p41_add_66886[16:3]};
  assign p42_add_68119_comb = {p41_add_67946[16:7] ^ p41_add_67946[18:9], p41_add_67946[6:0] ^ p41_add_67946[8:2] ^ p41_add_67946[31:25], p41_add_67946[31:30] ^ p41_add_67946[1:0] ^ p41_add_67946[24:23], p41_add_67946[29:17] ^ p41_add_67946[31:19] ^ p41_add_67946[22:10]} + p41_add_66752;
  assign p42_add_68022_comb = p42_add_68021_comb + p41_add_67551;
  assign p42_add_68028_comb = {p42_add_68025_comb, p41_add_67228[3:0]} + p41_add_67526;
  assign p42_add_68050_comb = p42_add_68048_comb + {p41_add_67893[1:0] ^ p41_add_67893[12:11] ^ p41_add_67893[21:20], p41_add_67893[31:21] ^ p41_add_67893[10:0] ^ p41_add_67893[19:9], p41_add_67893[20:12] ^ p41_add_67893[31:23] ^ p41_add_67893[8:0], p41_add_67893[11:2] ^ p41_add_67893[22:13] ^ p41_add_67893[31:22]};
  assign p42_add_68120_comb = p42_add_68118_comb + p42_add_68119_comb;
  assign p42_add_68137_comb = {p42_add_68085_comb[16:7] ^ p42_add_68085_comb[18:9], p42_add_68085_comb[6:0] ^ p42_add_68085_comb[8:2] ^ p42_add_68085_comb[31:25], p42_add_68085_comb[31:30] ^ p42_add_68085_comb[1:0] ^ p42_add_68085_comb[24:23], p42_add_68085_comb[29:17] ^ p42_add_68085_comb[31:19] ^ p42_add_68085_comb[22:10]} + p41_add_66886;
  assign p42_xor_68140_comb = p41_add_67228[3:0] ^ p41_add_67228[14:11] ^ p41_add_67228[31:28];

  // Registers for pipe stage 42:
  reg [31:0] p42_add_66921;
  reg [31:0] p42_add_67697;
  reg [31:0] p42_add_67059;
  reg [31:0] p42_add_67868;
  reg [31:0] p42_add_67094;
  reg [31:0] p42_add_68021;
  reg [31:0] p42_add_68022;
  reg [31:0] p42_add_67228;
  reg [31:0] p42_add_68028;
  reg [31:0] p42_add_67722;
  reg [31:0] p42_add_67263;
  reg [31:0] p42_add_67893;
  reg [31:0] p42_add_67400;
  reg [31:0] p42_and_68029;
  reg [31:0] p42_add_68050;
  reg [31:0] p42_add_67435;
  reg [1:0] p42_bit_slice_67552;
  reg [31:0] p42_add_67570;
  reg [31:0] p42_add_67604;
  reg [31:0] p42_add_67740;
  reg [31:0] p42_add_67775;
  reg [31:0] p42_add_67911;
  reg [1:0] p42_bit_slice_68051;
  reg [31:0] p42_add_67946;
  reg [31:0] p42_add_68085;
  reg [31:0] p42_add_68120;
  reg [31:0] p42_add_68137;
  reg [3:0] p42_xor_68140;
  always_ff @ (posedge clk) begin
    p42_add_66921 <= p41_add_66921;
    p42_add_67697 <= p41_add_67697;
    p42_add_67059 <= p41_add_67059;
    p42_add_67868 <= p41_add_67868;
    p42_add_67094 <= p41_add_67094;
    p42_add_68021 <= p42_add_68021_comb;
    p42_add_68022 <= p42_add_68022_comb;
    p42_add_67228 <= p41_add_67228;
    p42_add_68028 <= p42_add_68028_comb;
    p42_add_67722 <= p41_add_67722;
    p42_add_67263 <= p41_add_67263;
    p42_add_67893 <= p41_add_67893;
    p42_add_67400 <= p41_add_67400;
    p42_and_68029 <= p42_and_68029_comb;
    p42_add_68050 <= p42_add_68050_comb;
    p42_add_67435 <= p41_add_67435;
    p42_bit_slice_67552 <= p41_bit_slice_67552;
    p42_add_67570 <= p41_add_67570;
    p42_add_67604 <= p41_add_67604;
    p42_add_67740 <= p41_add_67740;
    p42_add_67775 <= p41_add_67775;
    p42_add_67911 <= p41_add_67911;
    p42_bit_slice_68051 <= p42_bit_slice_68051_comb;
    p42_add_67946 <= p41_add_67946;
    p42_add_68085 <= p42_add_68085_comb;
    p42_add_68120 <= p42_add_68120_comb;
    p42_add_68137 <= p42_add_68137_comb;
    p42_xor_68140 <= p42_xor_68140_comb;
  end

  // ===== Pipe stage 43:
  wire [31:0] p43_add_68262_comb;
  wire [31:0] p43_add_68263_comb;
  wire [31:0] p43_and_68224_comb;
  wire [31:0] p43_add_68218_comb;
  wire [31:0] p43_add_68219_comb;
  wire [31:0] p43_add_68222_comb;
  wire [31:0] p43_add_68243_comb;
  wire [31:0] p43_add_68296_comb;
  wire [31:0] p43_add_68297_comb;
  wire [31:0] p43_add_68220_comb;
  wire [31:0] p43_add_68223_comb;
  wire [31:0] p43_add_68245_comb;
  wire [31:0] p43_add_68298_comb;
  wire [31:0] p43_add_68315_comb;
  assign p43_add_68262_comb = p42_add_67604 + {p42_add_66921[6:4] ^ p42_add_66921[17:15], p42_add_66921[3:0] ^ p42_add_66921[14:11] ^ p42_add_66921[31:28], p42_add_66921[31:21] ^ p42_add_66921[10:0] ^ p42_add_66921[27:17], p42_add_66921[20:7] ^ p42_add_66921[31:18] ^ p42_add_66921[16:3]};
  assign p43_add_68263_comb = p43_add_68262_comb + p42_add_68137;
  assign p43_and_68224_comb = p42_add_68050 & p42_add_67893;
  assign p43_add_68218_comb = (p42_add_68022 & p42_add_67868 ^ ~(p42_add_68022 | ~p42_add_67697)) + {p42_add_68022[5:0] ^ p42_add_68022[10:5] ^ p42_add_68022[24:19], p42_add_68022[31:27] ^ p42_add_68022[4:0] ^ p42_add_68022[18:14], p42_add_68022[26:13] ^ p42_add_68022[31:18] ^ p42_add_68022[13:0], p42_add_68022[12:6] ^ p42_add_68022[17:11] ^ p42_add_68022[31:25]};
  assign p43_add_68219_comb = p43_add_68218_comb + p42_add_68028;
  assign p43_add_68222_comb = p42_add_67263 + 32'hc76c_51a3;
  assign p43_add_68243_comb = (p43_and_68224_comb ^ p42_add_68050 & p42_add_67722 ^ p42_and_68029) + p42_add_68021;
  assign p43_add_68296_comb = p42_add_67740 + {p42_add_67059[6:4] ^ p42_add_67059[17:15], p42_add_67059[3:0] ^ p42_add_67059[14:11] ^ p42_add_67059[31:28], p42_add_67059[31:21] ^ p42_add_67059[10:0] ^ p42_add_67059[27:17], p42_add_67059[20:7] ^ p42_add_67059[31:18] ^ p42_add_67059[16:3]};
  assign p43_add_68297_comb = {p42_add_68120[16:7] ^ p42_add_68120[18:9], p42_add_68120[6:0] ^ p42_add_68120[8:2] ^ p42_add_68120[31:25], p42_add_68120[31:30] ^ p42_add_68120[1:0] ^ p42_add_68120[24:23], p42_add_68120[29:17] ^ p42_add_68120[31:19] ^ p42_add_68120[22:10]} + p42_add_66921;
  assign p43_add_68220_comb = p43_add_68219_comb + p42_add_67722;
  assign p43_add_68223_comb = p42_add_67697 + p43_add_68222_comb;
  assign p43_add_68245_comb = p43_add_68243_comb + {p42_add_68050[1:0] ^ p42_add_68050[12:11] ^ p42_add_68050[21:20], p42_add_68050[31:21] ^ p42_add_68050[10:0] ^ p42_add_68050[19:9], p42_add_68050[20:12] ^ p42_add_68050[31:23] ^ p42_add_68050[8:0], p42_add_68050[11:2] ^ p42_add_68050[22:13] ^ p42_add_68050[31:22]};
  assign p43_add_68298_comb = p43_add_68296_comb + p43_add_68297_comb;
  assign p43_add_68315_comb = {p43_add_68263_comb[16:7] ^ p43_add_68263_comb[18:9], p43_add_68263_comb[6:0] ^ p43_add_68263_comb[8:2] ^ p43_add_68263_comb[31:25], p43_add_68263_comb[31:30] ^ p43_add_68263_comb[1:0] ^ p43_add_68263_comb[24:23], p43_add_68263_comb[29:17] ^ p43_add_68263_comb[31:19] ^ p43_add_68263_comb[22:10]} + p42_add_67059;

  // Registers for pipe stage 43:
  reg [31:0] p43_add_67868;
  reg [31:0] p43_add_67094;
  reg [31:0] p43_add_68022;
  reg [31:0] p43_add_67228;
  reg [31:0] p43_add_68219;
  reg [31:0] p43_add_68220;
  reg [31:0] p43_add_67263;
  reg [31:0] p43_add_68223;
  reg [31:0] p43_add_67893;
  reg [31:0] p43_add_67400;
  reg [31:0] p43_add_68050;
  reg [31:0] p43_add_67435;
  reg [1:0] p43_bit_slice_67552;
  reg [31:0] p43_and_68224;
  reg [31:0] p43_add_68245;
  reg [31:0] p43_add_67570;
  reg [31:0] p43_add_67604;
  reg [31:0] p43_add_67740;
  reg [31:0] p43_add_67775;
  reg [31:0] p43_add_67911;
  reg [1:0] p43_bit_slice_68051;
  reg [31:0] p43_add_67946;
  reg [31:0] p43_add_68085;
  reg [31:0] p43_add_68120;
  reg [31:0] p43_add_68263;
  reg [31:0] p43_add_68298;
  reg [31:0] p43_add_68315;
  reg [3:0] p43_xor_68140;
  always_ff @ (posedge clk) begin
    p43_add_67868 <= p42_add_67868;
    p43_add_67094 <= p42_add_67094;
    p43_add_68022 <= p42_add_68022;
    p43_add_67228 <= p42_add_67228;
    p43_add_68219 <= p43_add_68219_comb;
    p43_add_68220 <= p43_add_68220_comb;
    p43_add_67263 <= p42_add_67263;
    p43_add_68223 <= p43_add_68223_comb;
    p43_add_67893 <= p42_add_67893;
    p43_add_67400 <= p42_add_67400;
    p43_add_68050 <= p42_add_68050;
    p43_add_67435 <= p42_add_67435;
    p43_bit_slice_67552 <= p42_bit_slice_67552;
    p43_and_68224 <= p43_and_68224_comb;
    p43_add_68245 <= p43_add_68245_comb;
    p43_add_67570 <= p42_add_67570;
    p43_add_67604 <= p42_add_67604;
    p43_add_67740 <= p42_add_67740;
    p43_add_67775 <= p42_add_67775;
    p43_add_67911 <= p42_add_67911;
    p43_bit_slice_68051 <= p42_bit_slice_68051;
    p43_add_67946 <= p42_add_67946;
    p43_add_68085 <= p42_add_68085;
    p43_add_68120 <= p42_add_68120;
    p43_add_68263 <= p43_add_68263_comb;
    p43_add_68298 <= p43_add_68298_comb;
    p43_add_68315 <= p43_add_68315_comb;
    p43_xor_68140 <= p42_xor_68140;
  end

  // ===== Pipe stage 44:
  wire [31:0] p44_add_68446_comb;
  wire [31:0] p44_add_68447_comb;
  wire [31:0] p44_and_68399_comb;
  wire [31:0] p44_add_68393_comb;
  wire [31:0] p44_add_68394_comb;
  wire [31:0] p44_add_68397_comb;
  wire [31:0] p44_add_68418_comb;
  wire [28:0] p44_add_68423_comb;
  wire [29:0] p44_add_68428_comb;
  wire [31:0] p44_add_68476_comb;
  wire [31:0] p44_add_68477_comb;
  wire [31:0] p44_add_68395_comb;
  wire [31:0] p44_add_68398_comb;
  wire [31:0] p44_add_68420_comb;
  wire [31:0] p44_concat_68425_comb;
  wire [31:0] p44_concat_68429_comb;
  wire [31:0] p44_add_68478_comb;
  wire [31:0] p44_add_68495_comb;
  assign p44_add_68446_comb = p43_add_67775 + {p43_add_67094[6:4] ^ p43_add_67094[17:15], p43_add_67094[3:0] ^ p43_add_67094[14:11] ^ p43_add_67094[31:28], p43_add_67094[31:21] ^ p43_add_67094[10:0] ^ p43_add_67094[27:17], p43_add_67094[20:7] ^ p43_add_67094[31:18] ^ p43_add_67094[16:3]};
  assign p44_add_68447_comb = p44_add_68446_comb + p43_add_68315;
  assign p44_and_68399_comb = p43_add_68245 & p43_add_68050;
  assign p44_add_68393_comb = {p43_add_68220[5:0] ^ p43_add_68220[10:5] ^ p43_add_68220[24:19], p43_add_68220[31:27] ^ p43_add_68220[4:0] ^ p43_add_68220[18:14], p43_add_68220[26:13] ^ p43_add_68220[31:18] ^ p43_add_68220[13:0], p43_add_68220[12:6] ^ p43_add_68220[17:11] ^ p43_add_68220[31:25]} + (p43_add_68220 & p43_add_68022 ^ ~(p43_add_68220 | ~p43_add_67868));
  assign p44_add_68394_comb = p44_add_68393_comb + p43_add_68223;
  assign p44_add_68397_comb = p43_add_67400 + 32'hd192_e819;
  assign p44_add_68418_comb = (p44_and_68399_comb ^ p43_add_68245 & p43_add_67893 ^ p43_and_68224) + p43_add_68219;
  assign p44_add_68423_comb = p43_add_67775[31:3] + 29'h03c6_ed81;
  assign p44_add_68428_comb = p43_add_67911[31:2] + 30'h09d2_1dd3;
  assign p44_add_68476_comb = p43_add_67911 + {p43_add_67228[6:4] ^ p43_add_67228[17:15], p43_xor_68140, p43_add_67228[31:21] ^ p43_add_67228[10:0] ^ p43_add_67228[27:17], p43_add_67228[20:7] ^ p43_add_67228[31:18] ^ p43_add_67228[16:3]};
  assign p44_add_68477_comb = {p43_add_68298[16:7] ^ p43_add_68298[18:9], p43_add_68298[6:0] ^ p43_add_68298[8:2] ^ p43_add_68298[31:25], p43_add_68298[31:30] ^ p43_add_68298[1:0] ^ p43_add_68298[24:23], p43_add_68298[29:17] ^ p43_add_68298[31:19] ^ p43_add_68298[22:10]} + p43_add_67094;
  assign p44_add_68395_comb = p44_add_68394_comb + p43_add_67893;
  assign p44_add_68398_comb = p43_add_67868 + p44_add_68397_comb;
  assign p44_add_68420_comb = p44_add_68418_comb + {p43_add_68245[1:0] ^ p43_add_68245[12:11] ^ p43_add_68245[21:20], p43_add_68245[31:21] ^ p43_add_68245[10:0] ^ p43_add_68245[19:9], p43_add_68245[20:12] ^ p43_add_68245[31:23] ^ p43_add_68245[8:0], p43_add_68245[11:2] ^ p43_add_68245[22:13] ^ p43_add_68245[31:22]};
  assign p44_concat_68425_comb = {p44_add_68423_comb, p43_add_67775[2:0]};
  assign p44_concat_68429_comb = {p44_add_68428_comb, p43_bit_slice_68051};
  assign p44_add_68478_comb = p44_add_68476_comb + p44_add_68477_comb;
  assign p44_add_68495_comb = {p44_add_68447_comb[16:7] ^ p44_add_68447_comb[18:9], p44_add_68447_comb[6:0] ^ p44_add_68447_comb[8:2] ^ p44_add_68447_comb[31:25], p44_add_68447_comb[31:30] ^ p44_add_68447_comb[1:0] ^ p44_add_68447_comb[24:23], p44_add_68447_comb[29:17] ^ p44_add_68447_comb[31:19] ^ p44_add_68447_comb[22:10]} + p43_add_67228;

  // Registers for pipe stage 44:
  reg [31:0] p44_add_68022;
  reg [31:0] p44_add_68220;
  reg [31:0] p44_add_67263;
  reg [31:0] p44_add_68394;
  reg [31:0] p44_add_68395;
  reg [31:0] p44_add_67400;
  reg [31:0] p44_add_68398;
  reg [31:0] p44_add_68050;
  reg [31:0] p44_add_67435;
  reg [1:0] p44_bit_slice_67552;
  reg [31:0] p44_add_68245;
  reg [31:0] p44_add_67570;
  reg [31:0] p44_and_68399;
  reg [31:0] p44_add_68420;
  reg [31:0] p44_add_67604;
  reg [31:0] p44_add_67740;
  reg [31:0] p44_concat_68425;
  reg [31:0] p44_concat_68429;
  reg [31:0] p44_add_67946;
  reg [31:0] p44_add_68085;
  reg [31:0] p44_add_68120;
  reg [31:0] p44_add_68263;
  reg [31:0] p44_add_68298;
  reg [31:0] p44_add_68447;
  reg [31:0] p44_add_68478;
  reg [31:0] p44_add_68495;
  always_ff @ (posedge clk) begin
    p44_add_68022 <= p43_add_68022;
    p44_add_68220 <= p43_add_68220;
    p44_add_67263 <= p43_add_67263;
    p44_add_68394 <= p44_add_68394_comb;
    p44_add_68395 <= p44_add_68395_comb;
    p44_add_67400 <= p43_add_67400;
    p44_add_68398 <= p44_add_68398_comb;
    p44_add_68050 <= p43_add_68050;
    p44_add_67435 <= p43_add_67435;
    p44_bit_slice_67552 <= p43_bit_slice_67552;
    p44_add_68245 <= p43_add_68245;
    p44_add_67570 <= p43_add_67570;
    p44_and_68399 <= p44_and_68399_comb;
    p44_add_68420 <= p44_add_68420_comb;
    p44_add_67604 <= p43_add_67604;
    p44_add_67740 <= p43_add_67740;
    p44_concat_68425 <= p44_concat_68425_comb;
    p44_concat_68429 <= p44_concat_68429_comb;
    p44_add_67946 <= p43_add_67946;
    p44_add_68085 <= p43_add_68085;
    p44_add_68120 <= p43_add_68120;
    p44_add_68263 <= p43_add_68263;
    p44_add_68298 <= p43_add_68298;
    p44_add_68447 <= p44_add_68447_comb;
    p44_add_68478 <= p44_add_68478_comb;
    p44_add_68495 <= p44_add_68495_comb;
  end

  // ===== Pipe stage 45:
  wire [31:0] p45_add_68621_comb;
  wire [31:0] p45_add_68622_comb;
  wire [31:0] p45_and_68577_comb;
  wire [31:0] p45_add_68569_comb;
  wire [29:0] p45_add_68574_comb;
  wire [31:0] p45_add_68570_comb;
  wire [31:0] p45_add_68596_comb;
  wire [29:0] p45_add_68625_comb;
  wire [31:0] p45_add_68660_comb;
  wire [31:0] p45_add_68661_comb;
  wire [31:0] p45_add_68571_comb;
  wire [31:0] p45_add_68576_comb;
  wire [31:0] p45_add_68598_comb;
  wire [31:0] p45_add_68600_comb;
  wire [31:0] p45_add_68602_comb;
  wire [31:0] p45_add_68615_comb;
  wire [31:0] p45_concat_68649_comb;
  wire [31:0] p45_add_68662_comb;
  wire [31:0] p45_add_68678_comb;
  assign p45_add_68621_comb = p44_add_67946 + {p44_add_67263[6:4] ^ p44_add_67263[17:15], p44_add_67263[3:0] ^ p44_add_67263[14:11] ^ p44_add_67263[31:28], p44_add_67263[31:21] ^ p44_add_67263[10:0] ^ p44_add_67263[27:17], p44_add_67263[20:7] ^ p44_add_67263[31:18] ^ p44_add_67263[16:3]};
  assign p45_add_68622_comb = p45_add_68621_comb + p44_add_68495;
  assign p45_and_68577_comb = p44_add_68420 & p44_add_68245;
  assign p45_add_68569_comb = {p44_add_68395[5:0] ^ p44_add_68395[10:5] ^ p44_add_68395[24:19], p44_add_68395[31:27] ^ p44_add_68395[4:0] ^ p44_add_68395[18:14], p44_add_68395[26:13] ^ p44_add_68395[31:18] ^ p44_add_68395[13:0], p44_add_68395[12:6] ^ p44_add_68395[17:11] ^ p44_add_68395[31:25]} + (p44_add_68395 & p44_add_68220 ^ ~(p44_add_68395 | ~p44_add_68022));
  assign p45_add_68574_comb = p44_add_67435[31:2] + 30'h35a6_4189;
  assign p45_add_68570_comb = p45_add_68569_comb + p44_add_68398;
  assign p45_add_68596_comb = (p45_and_68577_comb ^ p44_add_68420 & p44_add_68050 ^ p44_and_68399) + p44_add_68394;
  assign p45_add_68625_comb = p45_add_68622_comb[31:2] + 30'h2132_1e05;
  assign p45_add_68660_comb = p44_add_68085 + {p44_add_67400[6:4] ^ p44_add_67400[17:15], p44_add_67400[3:0] ^ p44_add_67400[14:11] ^ p44_add_67400[31:28], p44_add_67400[31:21] ^ p44_add_67400[10:0] ^ p44_add_67400[27:17], p44_add_67400[20:7] ^ p44_add_67400[31:18] ^ p44_add_67400[16:3]};
  assign p45_add_68661_comb = {p44_add_68478[16:7] ^ p44_add_68478[18:9], p44_add_68478[6:0] ^ p44_add_68478[8:2] ^ p44_add_68478[31:25], p44_add_68478[31:30] ^ p44_add_68478[1:0] ^ p44_add_68478[24:23], p44_add_68478[29:17] ^ p44_add_68478[31:19] ^ p44_add_68478[22:10]} + p44_add_67263;
  assign p45_add_68571_comb = p45_add_68570_comb + p44_add_68050;
  assign p45_add_68576_comb = {p45_add_68574_comb, p44_bit_slice_67552} + p44_add_68022;
  assign p45_add_68598_comb = p45_add_68596_comb + {p44_add_68420[1:0] ^ p44_add_68420[12:11] ^ p44_add_68420[21:20], p44_add_68420[31:21] ^ p44_add_68420[10:0] ^ p44_add_68420[19:9], p44_add_68420[20:12] ^ p44_add_68420[31:23] ^ p44_add_68420[8:0], p44_add_68420[11:2] ^ p44_add_68420[22:13] ^ p44_add_68420[31:22]};
  assign p45_add_68600_comb = p44_add_67946 + 32'h34b0_bcb5;
  assign p45_add_68602_comb = p44_add_68085 + 32'h391c_0cb3;
  assign p45_add_68615_comb = p44_add_68478 + 32'h78a5_636f;
  assign p45_concat_68649_comb = {p45_add_68625_comb, p45_add_68622_comb[1:0]};
  assign p45_add_68662_comb = p45_add_68660_comb + p45_add_68661_comb;
  assign p45_add_68678_comb = {p45_add_68622_comb[16:7] ^ p45_add_68622_comb[18:9], p45_add_68622_comb[6:0] ^ p45_add_68622_comb[8:2] ^ p45_add_68622_comb[31:25], p45_add_68622_comb[31:30] ^ p45_add_68622_comb[1:0] ^ p45_add_68622_comb[24:23], p45_add_68622_comb[29:17] ^ p45_add_68622_comb[31:19] ^ p45_add_68622_comb[22:10]} + p44_add_67400;

  // Registers for pipe stage 45:
  reg [31:0] p45_add_68220;
  reg [31:0] p45_add_68395;
  reg [31:0] p45_add_68570;
  reg [31:0] p45_add_68571;
  reg [31:0] p45_add_67435;
  reg [31:0] p45_add_68576;
  reg [31:0] p45_add_68245;
  reg [31:0] p45_add_67570;
  reg [31:0] p45_add_68420;
  reg [31:0] p45_add_67604;
  reg [31:0] p45_and_68577;
  reg [31:0] p45_add_68598;
  reg [31:0] p45_add_67740;
  reg [31:0] p45_concat_68425;
  reg [31:0] p45_concat_68429;
  reg [31:0] p45_add_68600;
  reg [31:0] p45_add_68602;
  reg [31:0] p45_add_68120;
  reg [31:0] p45_add_68263;
  reg [31:0] p45_add_68298;
  reg [31:0] p45_add_68447;
  reg [31:0] p45_add_68615;
  reg [31:0] p45_concat_68649;
  reg [31:0] p45_add_68662;
  reg [31:0] p45_add_68678;
  always_ff @ (posedge clk) begin
    p45_add_68220 <= p44_add_68220;
    p45_add_68395 <= p44_add_68395;
    p45_add_68570 <= p45_add_68570_comb;
    p45_add_68571 <= p45_add_68571_comb;
    p45_add_67435 <= p44_add_67435;
    p45_add_68576 <= p45_add_68576_comb;
    p45_add_68245 <= p44_add_68245;
    p45_add_67570 <= p44_add_67570;
    p45_add_68420 <= p44_add_68420;
    p45_add_67604 <= p44_add_67604;
    p45_and_68577 <= p45_and_68577_comb;
    p45_add_68598 <= p45_add_68598_comb;
    p45_add_67740 <= p44_add_67740;
    p45_concat_68425 <= p44_concat_68425;
    p45_concat_68429 <= p44_concat_68429;
    p45_add_68600 <= p45_add_68600_comb;
    p45_add_68602 <= p45_add_68602_comb;
    p45_add_68120 <= p44_add_68120;
    p45_add_68263 <= p44_add_68263;
    p45_add_68298 <= p44_add_68298;
    p45_add_68447 <= p44_add_68447;
    p45_add_68615 <= p45_add_68615_comb;
    p45_concat_68649 <= p45_concat_68649_comb;
    p45_add_68662 <= p45_add_68662_comb;
    p45_add_68678 <= p45_add_68678_comb;
  end

  // ===== Pipe stage 46:
  wire [31:0] p46_and_68756_comb;
  wire [31:0] p46_add_68750_comb;
  wire [31:0] p46_add_68751_comb;
  wire [31:0] p46_add_68754_comb;
  wire [31:0] p46_add_68775_comb;
  wire [30:0] p46_add_68780_comb;
  wire [28:0] p46_add_68787_comb;
  wire [31:0] p46_add_68806_comb;
  wire [31:0] p46_add_68840_comb;
  wire [31:0] p46_add_68841_comb;
  wire [31:0] p46_add_68752_comb;
  wire [31:0] p46_add_68755_comb;
  wire [31:0] p46_add_68777_comb;
  wire [31:0] p46_concat_68782_comb;
  wire [31:0] p46_add_68784_comb;
  wire [31:0] p46_concat_68800_comb;
  wire [31:0] p46_add_68807_comb;
  wire [31:0] p46_add_68842_comb;
  assign p46_and_68756_comb = p45_add_68598 & p45_add_68420;
  assign p46_add_68750_comb = (p45_add_68571 & p45_add_68395 ^ ~(p45_add_68571 | ~p45_add_68220)) + {p45_add_68571[5:0] ^ p45_add_68571[10:5] ^ p45_add_68571[24:19], p45_add_68571[31:27] ^ p45_add_68571[4:0] ^ p45_add_68571[18:14], p45_add_68571[26:13] ^ p45_add_68571[31:18] ^ p45_add_68571[13:0], p45_add_68571[12:6] ^ p45_add_68571[17:11] ^ p45_add_68571[31:25]};
  assign p46_add_68751_comb = p46_add_68750_comb + p45_add_68576;
  assign p46_add_68754_comb = p45_add_67570 + 32'hf40e_3585;
  assign p46_add_68775_comb = (p46_and_68756_comb ^ p45_add_68598 & p45_add_68245 ^ p45_and_68577) + p45_add_68570;
  assign p46_add_68780_comb = p45_add_68120[31:1] + 31'h276c_5525;
  assign p46_add_68787_comb = p45_add_68662[31:3] + 29'h1198_e041;
  assign p46_add_68806_comb = p45_add_68120 + {p45_add_67435[6:4] ^ p45_add_67435[17:15], p45_add_67435[3:0] ^ p45_add_67435[14:11] ^ p45_add_67435[31:28], p45_add_67435[31:21] ^ p45_add_67435[10:0] ^ p45_add_67435[27:17], p45_add_67435[20:7] ^ p45_add_67435[31:18] ^ p45_add_67435[16:3]};
  assign p46_add_68840_comb = p45_add_68263 + {p45_add_67570[6:4] ^ p45_add_67570[17:15], p45_add_67570[3:0] ^ p45_add_67570[14:11] ^ p45_add_67570[31:28], p45_add_67570[31:21] ^ p45_add_67570[10:0] ^ p45_add_67570[27:17], p45_add_67570[20:7] ^ p45_add_67570[31:18] ^ p45_add_67570[16:3]};
  assign p46_add_68841_comb = {p45_add_68662[16:7] ^ p45_add_68662[18:9], p45_add_68662[6:0] ^ p45_add_68662[8:2] ^ p45_add_68662[31:25], p45_add_68662[31:30] ^ p45_add_68662[1:0] ^ p45_add_68662[24:23], p45_add_68662[29:17] ^ p45_add_68662[31:19] ^ p45_add_68662[22:10]} + p45_add_67435;
  assign p46_add_68752_comb = p46_add_68751_comb + p45_add_68245;
  assign p46_add_68755_comb = p45_add_68220 + p46_add_68754_comb;
  assign p46_add_68777_comb = p46_add_68775_comb + {p45_add_68598[1:0] ^ p45_add_68598[12:11] ^ p45_add_68598[21:20], p45_add_68598[31:21] ^ p45_add_68598[10:0] ^ p45_add_68598[19:9], p45_add_68598[20:12] ^ p45_add_68598[31:23] ^ p45_add_68598[8:0], p45_add_68598[11:2] ^ p45_add_68598[22:13] ^ p45_add_68598[31:22]};
  assign p46_concat_68782_comb = {p46_add_68780_comb, p45_add_68120[0]};
  assign p46_add_68784_comb = p45_add_68263 + 32'h5b9c_ca4f;
  assign p46_concat_68800_comb = {p46_add_68787_comb, p45_add_68662[2:0]};
  assign p46_add_68807_comb = p46_add_68806_comb + p45_add_68678;
  assign p46_add_68842_comb = p46_add_68840_comb + p46_add_68841_comb;

  // Registers for pipe stage 46:
  reg [31:0] p46_add_68395;
  reg [31:0] p46_add_68571;
  reg [31:0] p46_add_68751;
  reg [31:0] p46_add_68752;
  reg [31:0] p46_add_67570;
  reg [31:0] p46_add_68755;
  reg [31:0] p46_add_68420;
  reg [31:0] p46_add_67604;
  reg [31:0] p46_add_68598;
  reg [31:0] p46_add_67740;
  reg [31:0] p46_and_68756;
  reg [31:0] p46_add_68777;
  reg [31:0] p46_concat_68425;
  reg [31:0] p46_concat_68429;
  reg [31:0] p46_add_68600;
  reg [31:0] p46_add_68602;
  reg [31:0] p46_concat_68782;
  reg [31:0] p46_add_68784;
  reg [31:0] p46_add_68298;
  reg [31:0] p46_add_68447;
  reg [31:0] p46_add_68615;
  reg [31:0] p46_concat_68649;
  reg [31:0] p46_concat_68800;
  reg [31:0] p46_add_68807;
  reg [31:0] p46_add_68842;
  always_ff @ (posedge clk) begin
    p46_add_68395 <= p45_add_68395;
    p46_add_68571 <= p45_add_68571;
    p46_add_68751 <= p46_add_68751_comb;
    p46_add_68752 <= p46_add_68752_comb;
    p46_add_67570 <= p45_add_67570;
    p46_add_68755 <= p46_add_68755_comb;
    p46_add_68420 <= p45_add_68420;
    p46_add_67604 <= p45_add_67604;
    p46_add_68598 <= p45_add_68598;
    p46_add_67740 <= p45_add_67740;
    p46_and_68756 <= p46_and_68756_comb;
    p46_add_68777 <= p46_add_68777_comb;
    p46_concat_68425 <= p45_concat_68425;
    p46_concat_68429 <= p45_concat_68429;
    p46_add_68600 <= p45_add_68600;
    p46_add_68602 <= p45_add_68602;
    p46_concat_68782 <= p46_concat_68782_comb;
    p46_add_68784 <= p46_add_68784_comb;
    p46_add_68298 <= p45_add_68298;
    p46_add_68447 <= p45_add_68447;
    p46_add_68615 <= p45_add_68615;
    p46_concat_68649 <= p45_concat_68649;
    p46_concat_68800 <= p46_concat_68800_comb;
    p46_add_68807 <= p46_add_68807_comb;
    p46_add_68842 <= p46_add_68842_comb;
  end

  // ===== Pipe stage 47:
  wire [31:0] p47_and_68923_comb;
  wire [31:0] p47_add_68914_comb;
  wire [27:0] p47_add_68919_comb;
  wire [31:0] p47_add_68915_comb;
  wire [31:0] p47_add_68943_comb;
  wire [31:0] p47_add_68916_comb;
  wire [31:0] p47_add_68922_comb;
  wire [31:0] p47_add_68942_comb;
  wire [31:0] p47_add_68945_comb;
  wire [3:0] p47_xor_68948_comb;
  assign p47_and_68923_comb = p46_add_68777 & p46_add_68598;
  assign p47_add_68914_comb = {p46_add_68752[5:0] ^ p46_add_68752[10:5] ^ p46_add_68752[24:19], p46_add_68752[31:27] ^ p46_add_68752[4:0] ^ p46_add_68752[18:14], p46_add_68752[26:13] ^ p46_add_68752[31:18] ^ p46_add_68752[13:0], p46_add_68752[12:6] ^ p46_add_68752[17:11] ^ p46_add_68752[31:25]} + (p46_add_68752 & p46_add_68571 ^ ~(p46_add_68752 | ~p46_add_68395));
  assign p47_add_68919_comb = p46_add_67604[31:4] + 28'h106_aa07;
  assign p47_add_68915_comb = p47_add_68914_comb + p46_add_68755;
  assign p47_add_68943_comb = (p47_and_68923_comb ^ p46_add_68777 & p46_add_68420 ^ p46_and_68756) + p46_add_68751;
  assign p47_add_68916_comb = p47_add_68915_comb + p46_add_68420;
  assign p47_add_68922_comb = {p47_add_68919_comb, p46_add_67604[3:0]} + p46_add_68395;
  assign p47_add_68942_comb = p46_concat_68425 + p46_add_68752;
  assign p47_add_68945_comb = p47_add_68943_comb + {p46_add_68777[1:0] ^ p46_add_68777[12:11] ^ p46_add_68777[21:20], p46_add_68777[31:21] ^ p46_add_68777[10:0] ^ p46_add_68777[19:9], p46_add_68777[20:12] ^ p46_add_68777[31:23] ^ p46_add_68777[8:0], p46_add_68777[11:2] ^ p46_add_68777[22:13] ^ p46_add_68777[31:22]};
  assign p47_xor_68948_comb = p46_add_67604[3:0] ^ p46_add_67604[14:11] ^ p46_add_67604[31:28];

  // Registers for pipe stage 47:
  reg [31:0] p47_add_68571;
  reg [31:0] p47_add_68752;
  reg [31:0] p47_add_67570;
  reg [31:0] p47_add_68915;
  reg [31:0] p47_add_68916;
  reg [31:0] p47_add_67604;
  reg [31:0] p47_add_68922;
  reg [31:0] p47_add_68598;
  reg [31:0] p47_add_67740;
  reg [31:0] p47_add_68777;
  reg [31:0] p47_and_68923;
  reg [31:0] p47_add_68942;
  reg [31:0] p47_add_68945;
  reg [31:0] p47_concat_68429;
  reg [31:0] p47_add_68600;
  reg [31:0] p47_add_68602;
  reg [31:0] p47_concat_68782;
  reg [31:0] p47_add_68784;
  reg [31:0] p47_add_68298;
  reg [31:0] p47_add_68447;
  reg [31:0] p47_add_68615;
  reg [31:0] p47_concat_68649;
  reg [31:0] p47_concat_68800;
  reg [31:0] p47_add_68807;
  reg [31:0] p47_add_68842;
  reg [3:0] p47_xor_68948;
  always_ff @ (posedge clk) begin
    p47_add_68571 <= p46_add_68571;
    p47_add_68752 <= p46_add_68752;
    p47_add_67570 <= p46_add_67570;
    p47_add_68915 <= p47_add_68915_comb;
    p47_add_68916 <= p47_add_68916_comb;
    p47_add_67604 <= p46_add_67604;
    p47_add_68922 <= p47_add_68922_comb;
    p47_add_68598 <= p46_add_68598;
    p47_add_67740 <= p46_add_67740;
    p47_add_68777 <= p46_add_68777;
    p47_and_68923 <= p47_and_68923_comb;
    p47_add_68942 <= p47_add_68942_comb;
    p47_add_68945 <= p47_add_68945_comb;
    p47_concat_68429 <= p46_concat_68429;
    p47_add_68600 <= p46_add_68600;
    p47_add_68602 <= p46_add_68602;
    p47_concat_68782 <= p46_concat_68782;
    p47_add_68784 <= p46_add_68784;
    p47_add_68298 <= p46_add_68298;
    p47_add_68447 <= p46_add_68447;
    p47_add_68615 <= p46_add_68615;
    p47_concat_68649 <= p46_concat_68649;
    p47_concat_68800 <= p46_concat_68800;
    p47_add_68807 <= p46_add_68807;
    p47_add_68842 <= p46_add_68842;
    p47_xor_68948 <= p47_xor_68948_comb;
  end

  // ===== Pipe stage 48:
  wire [12:0] p48_xor_69074_comb;
  wire [31:0] p48_add_69022_comb;
  wire [31:0] p48_and_69033_comb;
  wire [31:0] p48_add_69023_comb;
  wire [30:0] p48_add_69029_comb;
  wire [30:0] p48_add_69097_comb;
  wire [31:0] p48_add_69024_comb;
  wire [31:0] p48_add_69053_comb;
  wire [30:0] p48_add_69058_comb;
  wire [31:0] p48_add_69099_comb;
  wire [31:0] p48_nor_69028_comb;
  wire [31:0] p48_add_69032_comb;
  wire [31:0] p48_add_69052_comb;
  wire [31:0] p48_add_69055_comb;
  wire [31:0] p48_concat_69060_comb;
  wire [31:0] p48_add_69062_comb;
  wire [31:0] p48_add_69101_comb;
  assign p48_xor_69074_comb = p47_add_68842[29:17] ^ p47_add_68842[31:19] ^ p47_add_68842[22:10];
  assign p48_add_69022_comb = (p47_add_68916 & p47_add_68752 ^ ~(p47_add_68916 | ~p47_add_68571)) + {p47_add_68916[5:0] ^ p47_add_68916[10:5] ^ p47_add_68916[24:19], p47_add_68916[31:27] ^ p47_add_68916[4:0] ^ p47_add_68916[18:14], p47_add_68916[26:13] ^ p47_add_68916[31:18] ^ p47_add_68916[13:0], p47_add_68916[12:6] ^ p47_add_68916[17:11] ^ p47_add_68916[31:25]};
  assign p48_and_69033_comb = p47_add_68945 & p47_add_68777;
  assign p48_add_69023_comb = p48_add_69022_comb + p47_add_68922;
  assign p48_add_69029_comb = p47_add_67740[31:1] + 31'h0cd2_608b;
  assign p48_add_69097_comb = {p47_add_68842[16:7] ^ p47_add_68842[18:9], p47_add_68842[6:0] ^ p47_add_68842[8:2] ^ p47_add_68842[31:25], p47_add_68842[31:30] ^ p47_add_68842[1:0] ^ p47_add_68842[24:23], p48_xor_69074_comb[12:1]} + 31'h6338_bc79;
  assign p48_add_69024_comb = p48_add_69023_comb + p47_add_68598;
  assign p48_add_69053_comb = (p48_and_69033_comb ^ p47_add_68945 & p47_add_68598 ^ p47_and_68923) + p47_add_68915;
  assign p48_add_69058_comb = p47_add_68447[31:1] + 31'h3a47_c177;
  assign p48_add_69099_comb = {p47_add_67740[6:4] ^ p47_add_67740[17:15], p47_add_67740[3:0] ^ p47_add_67740[14:11] ^ p47_add_67740[31:28], p47_add_67740[31:21] ^ p47_add_67740[10:0] ^ p47_add_67740[27:17], p47_add_67740[20:7] ^ p47_add_67740[31:18] ^ p47_add_67740[16:3]} + p47_add_68447;
  assign p48_nor_69028_comb = ~(p48_add_69024_comb | ~p47_add_68752);
  assign p48_add_69032_comb = {p48_add_69029_comb, p47_add_67740[0]} + p47_add_68571;
  assign p48_add_69052_comb = p47_concat_68429 + p47_add_68916;
  assign p48_add_69055_comb = p48_add_69053_comb + {p47_add_68945[1:0] ^ p47_add_68945[12:11] ^ p47_add_68945[21:20], p47_add_68945[31:21] ^ p47_add_68945[10:0] ^ p47_add_68945[19:9], p47_add_68945[20:12] ^ p47_add_68945[31:23] ^ p47_add_68945[8:0], p47_add_68945[11:2] ^ p47_add_68945[22:13] ^ p47_add_68945[31:22]};
  assign p48_concat_69060_comb = {p48_add_69058_comb, p47_add_68447[0]};
  assign p48_add_69062_comb = p47_add_68842 + 32'ha450_6ceb;
  assign p48_add_69101_comb = p48_add_69099_comb + {p48_add_69097_comb, p48_xor_69074_comb[0]};

  // Registers for pipe stage 48:
  reg [31:0] p48_add_67570;
  reg [31:0] p48_add_68916;
  reg [31:0] p48_add_67604;
  reg [31:0] p48_add_69023;
  reg [31:0] p48_add_69024;
  reg [31:0] p48_nor_69028;
  reg [31:0] p48_add_69032;
  reg [31:0] p48_add_68777;
  reg [31:0] p48_add_68942;
  reg [31:0] p48_add_68945;
  reg [31:0] p48_and_69033;
  reg [31:0] p48_add_69052;
  reg [31:0] p48_add_69055;
  reg [31:0] p48_add_68600;
  reg [31:0] p48_add_68602;
  reg [31:0] p48_concat_68782;
  reg [31:0] p48_add_68784;
  reg [31:0] p48_add_68298;
  reg [31:0] p48_concat_69060;
  reg [31:0] p48_add_68615;
  reg [31:0] p48_concat_68649;
  reg [31:0] p48_concat_68800;
  reg [31:0] p48_add_68807;
  reg [31:0] p48_add_69062;
  reg [3:0] p48_xor_68948;
  reg [31:0] p48_add_69101;
  always_ff @ (posedge clk) begin
    p48_add_67570 <= p47_add_67570;
    p48_add_68916 <= p47_add_68916;
    p48_add_67604 <= p47_add_67604;
    p48_add_69023 <= p48_add_69023_comb;
    p48_add_69024 <= p48_add_69024_comb;
    p48_nor_69028 <= p48_nor_69028_comb;
    p48_add_69032 <= p48_add_69032_comb;
    p48_add_68777 <= p47_add_68777;
    p48_add_68942 <= p47_add_68942;
    p48_add_68945 <= p47_add_68945;
    p48_and_69033 <= p48_and_69033_comb;
    p48_add_69052 <= p48_add_69052_comb;
    p48_add_69055 <= p48_add_69055_comb;
    p48_add_68600 <= p47_add_68600;
    p48_add_68602 <= p47_add_68602;
    p48_concat_68782 <= p47_concat_68782;
    p48_add_68784 <= p47_add_68784;
    p48_add_68298 <= p47_add_68298;
    p48_concat_69060 <= p48_concat_69060_comb;
    p48_add_68615 <= p47_add_68615;
    p48_concat_68649 <= p47_concat_68649;
    p48_concat_68800 <= p47_concat_68800;
    p48_add_68807 <= p47_add_68807;
    p48_add_69062 <= p48_add_69062_comb;
    p48_xor_68948 <= p47_xor_68948;
    p48_add_69101 <= p48_add_69101_comb;
  end

  // ===== Pipe stage 49:
  wire [31:0] p49_add_69173_comb;
  wire [31:0] p49_and_69178_comb;
  wire [31:0] p49_add_69174_comb;
  wire [31:0] p49_add_69175_comb;
  wire [31:0] p49_add_69198_comb;
  wire [31:0] p49_nor_69177_comb;
  wire [31:0] p49_add_69197_comb;
  wire [31:0] p49_add_69200_comb;
  assign p49_add_69173_comb = (p48_add_69024 & p48_add_68916 ^ p48_nor_69028) + {p48_add_69024[5:0] ^ p48_add_69024[10:5] ^ p48_add_69024[24:19], p48_add_69024[31:27] ^ p48_add_69024[4:0] ^ p48_add_69024[18:14], p48_add_69024[26:13] ^ p48_add_69024[31:18] ^ p48_add_69024[13:0], p48_add_69024[12:6] ^ p48_add_69024[17:11] ^ p48_add_69024[31:25]};
  assign p49_and_69178_comb = p48_add_69055 & p48_add_68945;
  assign p49_add_69174_comb = p49_add_69173_comb + p48_add_69032;
  assign p49_add_69175_comb = p49_add_69174_comb + p48_add_68777;
  assign p49_add_69198_comb = (p49_and_69178_comb ^ p48_add_69055 & p48_add_68777 ^ p48_and_69033) + p48_add_69023;
  assign p49_nor_69177_comb = ~(p49_add_69175_comb | ~p48_add_68916);
  assign p49_add_69197_comb = p48_add_69024 + p48_add_68600;
  assign p49_add_69200_comb = p49_add_69198_comb + {p48_add_69055[1:0] ^ p48_add_69055[12:11] ^ p48_add_69055[21:20], p48_add_69055[31:21] ^ p48_add_69055[10:0] ^ p48_add_69055[19:9], p48_add_69055[20:12] ^ p48_add_69055[31:23] ^ p48_add_69055[8:0], p48_add_69055[11:2] ^ p48_add_69055[22:13] ^ p48_add_69055[31:22]};

  // Registers for pipe stage 49:
  reg [31:0] p49_add_67570;
  reg [31:0] p49_add_67604;
  reg [31:0] p49_add_69024;
  reg [31:0] p49_add_69174;
  reg [31:0] p49_add_69175;
  reg [31:0] p49_nor_69177;
  reg [31:0] p49_add_68942;
  reg [31:0] p49_add_68945;
  reg [31:0] p49_add_69052;
  reg [31:0] p49_add_69055;
  reg [31:0] p49_and_69178;
  reg [31:0] p49_add_69197;
  reg [31:0] p49_add_69200;
  reg [31:0] p49_add_68602;
  reg [31:0] p49_concat_68782;
  reg [31:0] p49_add_68784;
  reg [31:0] p49_add_68298;
  reg [31:0] p49_concat_69060;
  reg [31:0] p49_add_68615;
  reg [31:0] p49_concat_68649;
  reg [31:0] p49_concat_68800;
  reg [31:0] p49_add_68807;
  reg [31:0] p49_add_69062;
  reg [3:0] p49_xor_68948;
  reg [31:0] p49_add_69101;
  always_ff @ (posedge clk) begin
    p49_add_67570 <= p48_add_67570;
    p49_add_67604 <= p48_add_67604;
    p49_add_69024 <= p48_add_69024;
    p49_add_69174 <= p49_add_69174_comb;
    p49_add_69175 <= p49_add_69175_comb;
    p49_nor_69177 <= p49_nor_69177_comb;
    p49_add_68942 <= p48_add_68942;
    p49_add_68945 <= p48_add_68945;
    p49_add_69052 <= p48_add_69052;
    p49_add_69055 <= p48_add_69055;
    p49_and_69178 <= p49_and_69178_comb;
    p49_add_69197 <= p49_add_69197_comb;
    p49_add_69200 <= p49_add_69200_comb;
    p49_add_68602 <= p48_add_68602;
    p49_concat_68782 <= p48_concat_68782;
    p49_add_68784 <= p48_add_68784;
    p49_add_68298 <= p48_add_68298;
    p49_concat_69060 <= p48_concat_69060;
    p49_add_68615 <= p48_add_68615;
    p49_concat_68649 <= p48_concat_68649;
    p49_concat_68800 <= p48_concat_68800;
    p49_add_68807 <= p48_add_68807;
    p49_add_69062 <= p48_add_69062;
    p49_xor_68948 <= p48_xor_68948;
    p49_add_69101 <= p48_add_69101;
  end

  // ===== Pipe stage 50:
  wire [31:0] p50_add_69270_comb;
  wire [31:0] p50_and_69275_comb;
  wire [31:0] p50_add_69271_comb;
  wire [31:0] p50_add_69272_comb;
  wire [31:0] p50_add_69295_comb;
  wire [31:0] p50_nor_69274_comb;
  wire [31:0] p50_add_69294_comb;
  wire [31:0] p50_add_69297_comb;
  assign p50_add_69270_comb = (p49_add_69175 & p49_add_69024 ^ p49_nor_69177) + {p49_add_69175[5:0] ^ p49_add_69175[10:5] ^ p49_add_69175[24:19], p49_add_69175[31:27] ^ p49_add_69175[4:0] ^ p49_add_69175[18:14], p49_add_69175[26:13] ^ p49_add_69175[31:18] ^ p49_add_69175[13:0], p49_add_69175[12:6] ^ p49_add_69175[17:11] ^ p49_add_69175[31:25]};
  assign p50_and_69275_comb = p49_add_69200 & p49_add_69055;
  assign p50_add_69271_comb = p50_add_69270_comb + p49_add_68942;
  assign p50_add_69272_comb = p50_add_69271_comb + p49_add_68945;
  assign p50_add_69295_comb = (p50_and_69275_comb ^ p49_add_69200 & p49_add_68945 ^ p49_and_69178) + p49_add_69174;
  assign p50_nor_69274_comb = ~(p50_add_69272_comb | ~p49_add_69024);
  assign p50_add_69294_comb = p49_add_69175 + p49_add_68602;
  assign p50_add_69297_comb = p50_add_69295_comb + {p49_add_69200[1:0] ^ p49_add_69200[12:11] ^ p49_add_69200[21:20], p49_add_69200[31:21] ^ p49_add_69200[10:0] ^ p49_add_69200[19:9], p49_add_69200[20:12] ^ p49_add_69200[31:23] ^ p49_add_69200[8:0], p49_add_69200[11:2] ^ p49_add_69200[22:13] ^ p49_add_69200[31:22]};

  // Registers for pipe stage 50:
  reg [31:0] p50_add_67570;
  reg [31:0] p50_add_67604;
  reg [31:0] p50_add_69175;
  reg [31:0] p50_add_69271;
  reg [31:0] p50_add_69272;
  reg [31:0] p50_nor_69274;
  reg [31:0] p50_add_69052;
  reg [31:0] p50_add_69055;
  reg [31:0] p50_add_69197;
  reg [31:0] p50_add_69200;
  reg [31:0] p50_and_69275;
  reg [31:0] p50_add_69294;
  reg [31:0] p50_add_69297;
  reg [31:0] p50_concat_68782;
  reg [31:0] p50_add_68784;
  reg [31:0] p50_add_68298;
  reg [31:0] p50_concat_69060;
  reg [31:0] p50_add_68615;
  reg [31:0] p50_concat_68649;
  reg [31:0] p50_concat_68800;
  reg [31:0] p50_add_68807;
  reg [31:0] p50_add_69062;
  reg [3:0] p50_xor_68948;
  reg [31:0] p50_add_69101;
  always_ff @ (posedge clk) begin
    p50_add_67570 <= p49_add_67570;
    p50_add_67604 <= p49_add_67604;
    p50_add_69175 <= p49_add_69175;
    p50_add_69271 <= p50_add_69271_comb;
    p50_add_69272 <= p50_add_69272_comb;
    p50_nor_69274 <= p50_nor_69274_comb;
    p50_add_69052 <= p49_add_69052;
    p50_add_69055 <= p49_add_69055;
    p50_add_69197 <= p49_add_69197;
    p50_add_69200 <= p49_add_69200;
    p50_and_69275 <= p50_and_69275_comb;
    p50_add_69294 <= p50_add_69294_comb;
    p50_add_69297 <= p50_add_69297_comb;
    p50_concat_68782 <= p49_concat_68782;
    p50_add_68784 <= p49_add_68784;
    p50_add_68298 <= p49_add_68298;
    p50_concat_69060 <= p49_concat_69060;
    p50_add_68615 <= p49_add_68615;
    p50_concat_68649 <= p49_concat_68649;
    p50_concat_68800 <= p49_concat_68800;
    p50_add_68807 <= p49_add_68807;
    p50_add_69062 <= p49_add_69062;
    p50_xor_68948 <= p49_xor_68948;
    p50_add_69101 <= p49_add_69101;
  end

  // ===== Pipe stage 51:
  wire [31:0] p51_add_69365_comb;
  wire [31:0] p51_and_69370_comb;
  wire [31:0] p51_add_69366_comb;
  wire [31:0] p51_add_69367_comb;
  wire [31:0] p51_add_69390_comb;
  wire [31:0] p51_nor_69369_comb;
  wire [31:0] p51_add_69389_comb;
  wire [31:0] p51_add_69392_comb;
  assign p51_add_69365_comb = (p50_add_69272 & p50_add_69175 ^ p50_nor_69274) + {p50_add_69272[5:0] ^ p50_add_69272[10:5] ^ p50_add_69272[24:19], p50_add_69272[31:27] ^ p50_add_69272[4:0] ^ p50_add_69272[18:14], p50_add_69272[26:13] ^ p50_add_69272[31:18] ^ p50_add_69272[13:0], p50_add_69272[12:6] ^ p50_add_69272[17:11] ^ p50_add_69272[31:25]};
  assign p51_and_69370_comb = p50_add_69297 & p50_add_69200;
  assign p51_add_69366_comb = p51_add_69365_comb + p50_add_69052;
  assign p51_add_69367_comb = p51_add_69366_comb + p50_add_69055;
  assign p51_add_69390_comb = (p51_and_69370_comb ^ p50_add_69297 & p50_add_69055 ^ p50_and_69275) + p50_add_69271;
  assign p51_nor_69369_comb = ~(p51_add_69367_comb | ~p50_add_69175);
  assign p51_add_69389_comb = p50_concat_68782 + p50_add_69272;
  assign p51_add_69392_comb = p51_add_69390_comb + {p50_add_69297[1:0] ^ p50_add_69297[12:11] ^ p50_add_69297[21:20], p50_add_69297[31:21] ^ p50_add_69297[10:0] ^ p50_add_69297[19:9], p50_add_69297[20:12] ^ p50_add_69297[31:23] ^ p50_add_69297[8:0], p50_add_69297[11:2] ^ p50_add_69297[22:13] ^ p50_add_69297[31:22]};

  // Registers for pipe stage 51:
  reg [31:0] p51_add_67570;
  reg [31:0] p51_add_67604;
  reg [31:0] p51_add_69272;
  reg [31:0] p51_add_69366;
  reg [31:0] p51_add_69367;
  reg [31:0] p51_nor_69369;
  reg [31:0] p51_add_69197;
  reg [31:0] p51_add_69200;
  reg [31:0] p51_add_69294;
  reg [31:0] p51_add_69297;
  reg [31:0] p51_and_69370;
  reg [31:0] p51_add_69389;
  reg [31:0] p51_add_69392;
  reg [31:0] p51_add_68784;
  reg [31:0] p51_add_68298;
  reg [31:0] p51_concat_69060;
  reg [31:0] p51_add_68615;
  reg [31:0] p51_concat_68649;
  reg [31:0] p51_concat_68800;
  reg [31:0] p51_add_68807;
  reg [31:0] p51_add_69062;
  reg [3:0] p51_xor_68948;
  reg [31:0] p51_add_69101;
  always_ff @ (posedge clk) begin
    p51_add_67570 <= p50_add_67570;
    p51_add_67604 <= p50_add_67604;
    p51_add_69272 <= p50_add_69272;
    p51_add_69366 <= p51_add_69366_comb;
    p51_add_69367 <= p51_add_69367_comb;
    p51_nor_69369 <= p51_nor_69369_comb;
    p51_add_69197 <= p50_add_69197;
    p51_add_69200 <= p50_add_69200;
    p51_add_69294 <= p50_add_69294;
    p51_add_69297 <= p50_add_69297;
    p51_and_69370 <= p51_and_69370_comb;
    p51_add_69389 <= p51_add_69389_comb;
    p51_add_69392 <= p51_add_69392_comb;
    p51_add_68784 <= p50_add_68784;
    p51_add_68298 <= p50_add_68298;
    p51_concat_69060 <= p50_concat_69060;
    p51_add_68615 <= p50_add_68615;
    p51_concat_68649 <= p50_concat_68649;
    p51_concat_68800 <= p50_concat_68800;
    p51_add_68807 <= p50_add_68807;
    p51_add_69062 <= p50_add_69062;
    p51_xor_68948 <= p50_xor_68948;
    p51_add_69101 <= p50_add_69101;
  end

  // ===== Pipe stage 52:
  wire [31:0] p52_add_69458_comb;
  wire [31:0] p52_and_69463_comb;
  wire [31:0] p52_add_69459_comb;
  wire [31:0] p52_add_69460_comb;
  wire [31:0] p52_add_69483_comb;
  wire [31:0] p52_nor_69462_comb;
  wire [31:0] p52_add_69482_comb;
  wire [31:0] p52_add_69485_comb;
  assign p52_add_69458_comb = {p51_add_69367[5:0] ^ p51_add_69367[10:5] ^ p51_add_69367[24:19], p51_add_69367[31:27] ^ p51_add_69367[4:0] ^ p51_add_69367[18:14], p51_add_69367[26:13] ^ p51_add_69367[31:18] ^ p51_add_69367[13:0], p51_add_69367[12:6] ^ p51_add_69367[17:11] ^ p51_add_69367[31:25]} + (p51_add_69367 & p51_add_69272 ^ p51_nor_69369);
  assign p52_and_69463_comb = p51_add_69392 & p51_add_69297;
  assign p52_add_69459_comb = p52_add_69458_comb + p51_add_69197;
  assign p52_add_69460_comb = p52_add_69459_comb + p51_add_69200;
  assign p52_add_69483_comb = (p52_and_69463_comb ^ p51_add_69392 & p51_add_69200 ^ p51_and_69370) + p51_add_69366;
  assign p52_nor_69462_comb = ~(p52_add_69460_comb | ~p51_add_69272);
  assign p52_add_69482_comb = p51_add_69367 + p51_add_68784;
  assign p52_add_69485_comb = p52_add_69483_comb + {p51_add_69392[1:0] ^ p51_add_69392[12:11] ^ p51_add_69392[21:20], p51_add_69392[31:21] ^ p51_add_69392[10:0] ^ p51_add_69392[19:9], p51_add_69392[20:12] ^ p51_add_69392[31:23] ^ p51_add_69392[8:0], p51_add_69392[11:2] ^ p51_add_69392[22:13] ^ p51_add_69392[31:22]};

  // Registers for pipe stage 52:
  reg [31:0] p52_add_67570;
  reg [31:0] p52_add_67604;
  reg [31:0] p52_add_69367;
  reg [31:0] p52_add_69459;
  reg [31:0] p52_add_69460;
  reg [31:0] p52_nor_69462;
  reg [31:0] p52_add_69294;
  reg [31:0] p52_add_69297;
  reg [31:0] p52_add_69389;
  reg [31:0] p52_add_69392;
  reg [31:0] p52_and_69463;
  reg [31:0] p52_add_69482;
  reg [31:0] p52_add_69485;
  reg [31:0] p52_add_68298;
  reg [31:0] p52_concat_69060;
  reg [31:0] p52_add_68615;
  reg [31:0] p52_concat_68649;
  reg [31:0] p52_concat_68800;
  reg [31:0] p52_add_68807;
  reg [31:0] p52_add_69062;
  reg [3:0] p52_xor_68948;
  reg [31:0] p52_add_69101;
  always_ff @ (posedge clk) begin
    p52_add_67570 <= p51_add_67570;
    p52_add_67604 <= p51_add_67604;
    p52_add_69367 <= p51_add_69367;
    p52_add_69459 <= p52_add_69459_comb;
    p52_add_69460 <= p52_add_69460_comb;
    p52_nor_69462 <= p52_nor_69462_comb;
    p52_add_69294 <= p51_add_69294;
    p52_add_69297 <= p51_add_69297;
    p52_add_69389 <= p51_add_69389;
    p52_add_69392 <= p51_add_69392;
    p52_and_69463 <= p52_and_69463_comb;
    p52_add_69482 <= p52_add_69482_comb;
    p52_add_69485 <= p52_add_69485_comb;
    p52_add_68298 <= p51_add_68298;
    p52_concat_69060 <= p51_concat_69060;
    p52_add_68615 <= p51_add_68615;
    p52_concat_68649 <= p51_concat_68649;
    p52_concat_68800 <= p51_concat_68800;
    p52_add_68807 <= p51_add_68807;
    p52_add_69062 <= p51_add_69062;
    p52_xor_68948 <= p51_xor_68948;
    p52_add_69101 <= p51_add_69101;
  end

  // ===== Pipe stage 53:
  wire [31:0] p53_add_69549_comb;
  wire [31:0] p53_and_69554_comb;
  wire [31:0] p53_add_69550_comb;
  wire [31:0] p53_add_69551_comb;
  wire [31:0] p53_add_69573_comb;
  wire [31:0] p53_nor_69553_comb;
  wire [31:0] p53_add_69575_comb;
  assign p53_add_69549_comb = {p52_add_69460[5:0] ^ p52_add_69460[10:5] ^ p52_add_69460[24:19], p52_add_69460[31:27] ^ p52_add_69460[4:0] ^ p52_add_69460[18:14], p52_add_69460[26:13] ^ p52_add_69460[31:18] ^ p52_add_69460[13:0], p52_add_69460[12:6] ^ p52_add_69460[17:11] ^ p52_add_69460[31:25]} + (p52_add_69460 & p52_add_69367 ^ p52_nor_69462);
  assign p53_and_69554_comb = p52_add_69485 & p52_add_69392;
  assign p53_add_69550_comb = p53_add_69549_comb + p52_add_69294;
  assign p53_add_69551_comb = p53_add_69550_comb + p52_add_69297;
  assign p53_add_69573_comb = (p53_and_69554_comb ^ p52_add_69485 & p52_add_69297 ^ p52_and_69463) + p52_add_69459;
  assign p53_nor_69553_comb = ~(p53_add_69551_comb | ~p52_add_69367);
  assign p53_add_69575_comb = p53_add_69573_comb + {p52_add_69485[1:0] ^ p52_add_69485[12:11] ^ p52_add_69485[21:20], p52_add_69485[31:21] ^ p52_add_69485[10:0] ^ p52_add_69485[19:9], p52_add_69485[20:12] ^ p52_add_69485[31:23] ^ p52_add_69485[8:0], p52_add_69485[11:2] ^ p52_add_69485[22:13] ^ p52_add_69485[31:22]};

  // Registers for pipe stage 53:
  reg [31:0] p53_add_67570;
  reg [31:0] p53_add_67604;
  reg [31:0] p53_add_69460;
  reg [31:0] p53_add_69550;
  reg [31:0] p53_add_69551;
  reg [31:0] p53_nor_69553;
  reg [31:0] p53_add_69389;
  reg [31:0] p53_add_69392;
  reg [31:0] p53_add_69482;
  reg [31:0] p53_add_69485;
  reg [31:0] p53_add_68298;
  reg [31:0] p53_and_69554;
  reg [31:0] p53_add_69575;
  reg [31:0] p53_concat_69060;
  reg [31:0] p53_add_68615;
  reg [31:0] p53_concat_68649;
  reg [31:0] p53_concat_68800;
  reg [31:0] p53_add_68807;
  reg [31:0] p53_add_69062;
  reg [3:0] p53_xor_68948;
  reg [31:0] p53_add_69101;
  always_ff @ (posedge clk) begin
    p53_add_67570 <= p52_add_67570;
    p53_add_67604 <= p52_add_67604;
    p53_add_69460 <= p52_add_69460;
    p53_add_69550 <= p53_add_69550_comb;
    p53_add_69551 <= p53_add_69551_comb;
    p53_nor_69553 <= p53_nor_69553_comb;
    p53_add_69389 <= p52_add_69389;
    p53_add_69392 <= p52_add_69392;
    p53_add_69482 <= p52_add_69482;
    p53_add_69485 <= p52_add_69485;
    p53_add_68298 <= p52_add_68298;
    p53_and_69554 <= p53_and_69554_comb;
    p53_add_69575 <= p53_add_69575_comb;
    p53_concat_69060 <= p52_concat_69060;
    p53_add_68615 <= p52_add_68615;
    p53_concat_68649 <= p52_concat_68649;
    p53_concat_68800 <= p52_concat_68800;
    p53_add_68807 <= p52_add_68807;
    p53_add_69062 <= p52_add_69062;
    p53_xor_68948 <= p52_xor_68948;
    p53_add_69101 <= p52_add_69101;
  end

  // ===== Pipe stage 54:
  wire [31:0] p54_and_69640_comb;
  wire [31:0] p54_add_69637_comb;
  wire [31:0] p54_add_69638_comb;
  wire [31:0] p54_add_69660_comb;
  wire [31:0] p54_add_69639_comb;
  wire [31:0] p54_add_69659_comb;
  wire [31:0] p54_add_69662_comb;
  assign p54_and_69640_comb = p53_add_69575 & p53_add_69485;
  assign p54_add_69637_comb = (p53_add_69551 & p53_add_69460 ^ p53_nor_69553) + {p53_add_69551[5:0] ^ p53_add_69551[10:5] ^ p53_add_69551[24:19], p53_add_69551[31:27] ^ p53_add_69551[4:0] ^ p53_add_69551[18:14], p53_add_69551[26:13] ^ p53_add_69551[31:18] ^ p53_add_69551[13:0], p53_add_69551[12:6] ^ p53_add_69551[17:11] ^ p53_add_69551[31:25]};
  assign p54_add_69638_comb = p54_add_69637_comb + p53_add_69389;
  assign p54_add_69660_comb = (p54_and_69640_comb ^ p53_add_69575 & p53_add_69392 ^ p53_and_69554) + p53_add_69550;
  assign p54_add_69639_comb = p54_add_69638_comb + p53_add_69392;
  assign p54_add_69659_comb = p53_concat_69060 + p53_add_69551;
  assign p54_add_69662_comb = p54_add_69660_comb + {p53_add_69575[1:0] ^ p53_add_69575[12:11] ^ p53_add_69575[21:20], p53_add_69575[31:21] ^ p53_add_69575[10:0] ^ p53_add_69575[19:9], p53_add_69575[20:12] ^ p53_add_69575[31:23] ^ p53_add_69575[8:0], p53_add_69575[11:2] ^ p53_add_69575[22:13] ^ p53_add_69575[31:22]};

  // Registers for pipe stage 54:
  reg [31:0] p54_add_67570;
  reg [31:0] p54_add_67604;
  reg [31:0] p54_add_69460;
  reg [31:0] p54_add_69551;
  reg [31:0] p54_add_69638;
  reg [31:0] p54_add_69639;
  reg [31:0] p54_add_69482;
  reg [31:0] p54_add_69485;
  reg [31:0] p54_add_68298;
  reg [31:0] p54_add_69575;
  reg [31:0] p54_and_69640;
  reg [31:0] p54_add_69659;
  reg [31:0] p54_add_69662;
  reg [31:0] p54_add_68615;
  reg [31:0] p54_concat_68649;
  reg [31:0] p54_concat_68800;
  reg [31:0] p54_add_68807;
  reg [31:0] p54_add_69062;
  reg [3:0] p54_xor_68948;
  reg [31:0] p54_add_69101;
  always_ff @ (posedge clk) begin
    p54_add_67570 <= p53_add_67570;
    p54_add_67604 <= p53_add_67604;
    p54_add_69460 <= p53_add_69460;
    p54_add_69551 <= p53_add_69551;
    p54_add_69638 <= p54_add_69638_comb;
    p54_add_69639 <= p54_add_69639_comb;
    p54_add_69482 <= p53_add_69482;
    p54_add_69485 <= p53_add_69485;
    p54_add_68298 <= p53_add_68298;
    p54_add_69575 <= p53_add_69575;
    p54_and_69640 <= p54_and_69640_comb;
    p54_add_69659 <= p54_add_69659_comb;
    p54_add_69662 <= p54_add_69662_comb;
    p54_add_68615 <= p53_add_68615;
    p54_concat_68649 <= p53_concat_68649;
    p54_concat_68800 <= p53_concat_68800;
    p54_add_68807 <= p53_add_68807;
    p54_add_69062 <= p53_add_69062;
    p54_xor_68948 <= p53_xor_68948;
    p54_add_69101 <= p53_add_69101;
  end

  // ===== Pipe stage 55:
  wire [31:0] p55_add_69724_comb;
  wire [31:0] p55_and_69732_comb;
  wire [31:0] p55_add_69725_comb;
  wire [31:0] p55_add_69726_comb;
  wire [31:0] p55_add_69730_comb;
  wire [31:0] p55_add_69751_comb;
  wire [30:0] p55_add_69757_comb;
  wire [31:0] p55_add_69789_comb;
  wire [31:0] p55_add_69790_comb;
  wire [31:0] p55_nor_69728_comb;
  wire [31:0] p55_add_69731_comb;
  wire [31:0] p55_add_69753_comb;
  wire [31:0] p55_add_69754_comb;
  wire [31:0] p55_concat_69759_comb;
  wire [31:0] p55_add_69791_comb;
  assign p55_add_69724_comb = {p54_add_69639[5:0] ^ p54_add_69639[10:5] ^ p54_add_69639[24:19], p54_add_69639[31:27] ^ p54_add_69639[4:0] ^ p54_add_69639[18:14], p54_add_69639[26:13] ^ p54_add_69639[31:18] ^ p54_add_69639[13:0], p54_add_69639[12:6] ^ p54_add_69639[17:11] ^ p54_add_69639[31:25]} + (p54_add_69639 & p54_add_69551 ^ ~(p54_add_69639 | ~p54_add_69460));
  assign p55_and_69732_comb = p54_add_69662 & p54_add_69575;
  assign p55_add_69725_comb = p55_add_69724_comb + p54_add_69482;
  assign p55_add_69726_comb = p55_add_69725_comb + p54_add_69485;
  assign p55_add_69730_comb = p54_add_68298 + 32'h682e_6ff3;
  assign p55_add_69751_comb = (p55_and_69732_comb ^ p54_add_69662 & p54_add_69485 ^ p54_and_69640) + p54_add_69638;
  assign p55_add_69757_comb = p54_add_68807[31:1] + 31'h485f_7ffd;
  assign p55_add_69789_comb = {p54_add_67604[6:4] ^ p54_add_67604[17:15], p54_xor_68948, p54_add_67604[31:21] ^ p54_add_67604[10:0] ^ p54_add_67604[27:17], p54_add_67604[20:7] ^ p54_add_67604[31:18] ^ p54_add_67604[16:3]} + p54_add_68298;
  assign p55_add_69790_comb = {p54_add_68807[16:7] ^ p54_add_68807[18:9], p54_add_68807[6:0] ^ p54_add_68807[8:2] ^ p54_add_68807[31:25], p54_add_68807[31:30] ^ p54_add_68807[1:0] ^ p54_add_68807[24:23], p54_add_68807[29:17] ^ p54_add_68807[31:19] ^ p54_add_68807[22:10]} + 32'hbef9_a3f7;
  assign p55_nor_69728_comb = ~(p55_add_69726_comb | ~p54_add_69551);
  assign p55_add_69731_comb = p54_add_69460 + p55_add_69730_comb;
  assign p55_add_69753_comb = p55_add_69751_comb + {p54_add_69662[1:0] ^ p54_add_69662[12:11] ^ p54_add_69662[21:20], p54_add_69662[31:21] ^ p54_add_69662[10:0] ^ p54_add_69662[19:9], p54_add_69662[20:12] ^ p54_add_69662[31:23] ^ p54_add_69662[8:0], p54_add_69662[11:2] ^ p54_add_69662[22:13] ^ p54_add_69662[31:22]};
  assign p55_add_69754_comb = p54_add_69639 + p54_add_68615;
  assign p55_concat_69759_comb = {p55_add_69757_comb, p54_add_68807[0]};
  assign p55_add_69791_comb = p55_add_69789_comb + p55_add_69790_comb;

  // Registers for pipe stage 55:
  reg [31:0] p55_add_67570;
  reg [31:0] p55_add_67604;
  reg [31:0] p55_add_69639;
  reg [31:0] p55_add_69725;
  reg [31:0] p55_add_69726;
  reg [31:0] p55_nor_69728;
  reg [31:0] p55_add_69731;
  reg [31:0] p55_add_69575;
  reg [31:0] p55_add_69659;
  reg [31:0] p55_add_69662;
  reg [31:0] p55_and_69732;
  reg [31:0] p55_add_69753;
  reg [31:0] p55_add_69754;
  reg [31:0] p55_concat_68649;
  reg [31:0] p55_concat_68800;
  reg [31:0] p55_concat_69759;
  reg [31:0] p55_add_69062;
  reg [31:0] p55_add_69101;
  reg [31:0] p55_add_69791;
  always_ff @ (posedge clk) begin
    p55_add_67570 <= p54_add_67570;
    p55_add_67604 <= p54_add_67604;
    p55_add_69639 <= p54_add_69639;
    p55_add_69725 <= p55_add_69725_comb;
    p55_add_69726 <= p55_add_69726_comb;
    p55_nor_69728 <= p55_nor_69728_comb;
    p55_add_69731 <= p55_add_69731_comb;
    p55_add_69575 <= p54_add_69575;
    p55_add_69659 <= p54_add_69659;
    p55_add_69662 <= p54_add_69662;
    p55_and_69732 <= p55_and_69732_comb;
    p55_add_69753 <= p55_add_69753_comb;
    p55_add_69754 <= p55_add_69754_comb;
    p55_concat_68649 <= p54_concat_68649;
    p55_concat_68800 <= p54_concat_68800;
    p55_concat_69759 <= p55_concat_69759_comb;
    p55_add_69062 <= p54_add_69062;
    p55_add_69101 <= p54_add_69101;
    p55_add_69791 <= p55_add_69791_comb;
  end

  // ===== Pipe stage 56:
  wire [31:0] p56_add_69849_comb;
  wire [31:0] p56_and_69854_comb;
  wire [31:0] p56_add_69850_comb;
  wire [31:0] p56_add_69851_comb;
  wire [31:0] p56_add_69873_comb;
  wire [31:0] p56_nor_69853_comb;
  wire [31:0] p56_add_69875_comb;
  wire [31:0] p56_add_69876_comb;
  assign p56_add_69849_comb = {p55_add_69726[5:0] ^ p55_add_69726[10:5] ^ p55_add_69726[24:19], p55_add_69726[31:27] ^ p55_add_69726[4:0] ^ p55_add_69726[18:14], p55_add_69726[26:13] ^ p55_add_69726[31:18] ^ p55_add_69726[13:0], p55_add_69726[12:6] ^ p55_add_69726[17:11] ^ p55_add_69726[31:25]} + (p55_add_69726 & p55_add_69639 ^ p55_nor_69728);
  assign p56_and_69854_comb = p55_add_69753 & p55_add_69662;
  assign p56_add_69850_comb = p56_add_69849_comb + p55_add_69731;
  assign p56_add_69851_comb = p56_add_69850_comb + p55_add_69575;
  assign p56_add_69873_comb = (p56_and_69854_comb ^ p55_add_69753 & p55_add_69575 ^ p55_and_69732) + p55_add_69725;
  assign p56_nor_69853_comb = ~(p56_add_69851_comb | ~p55_add_69639);
  assign p56_add_69875_comb = p56_add_69873_comb + {p55_add_69753[1:0] ^ p55_add_69753[12:11] ^ p55_add_69753[21:20], p55_add_69753[31:21] ^ p55_add_69753[10:0] ^ p55_add_69753[19:9], p55_add_69753[20:12] ^ p55_add_69753[31:23] ^ p55_add_69753[8:0], p55_add_69753[11:2] ^ p55_add_69753[22:13] ^ p55_add_69753[31:22]};
  assign p56_add_69876_comb = p55_concat_68649 + p55_add_69726;

  // Registers for pipe stage 56:
  reg [31:0] p56_add_67570;
  reg [31:0] p56_add_67604;
  reg [31:0] p56_add_69726;
  reg [31:0] p56_add_69850;
  reg [31:0] p56_add_69851;
  reg [31:0] p56_nor_69853;
  reg [31:0] p56_add_69659;
  reg [31:0] p56_add_69662;
  reg [31:0] p56_add_69753;
  reg [31:0] p56_add_69754;
  reg [31:0] p56_and_69854;
  reg [31:0] p56_add_69875;
  reg [31:0] p56_add_69876;
  reg [31:0] p56_concat_68800;
  reg [31:0] p56_concat_69759;
  reg [31:0] p56_add_69062;
  reg [31:0] p56_add_69101;
  reg [31:0] p56_add_69791;
  always_ff @ (posedge clk) begin
    p56_add_67570 <= p55_add_67570;
    p56_add_67604 <= p55_add_67604;
    p56_add_69726 <= p55_add_69726;
    p56_add_69850 <= p56_add_69850_comb;
    p56_add_69851 <= p56_add_69851_comb;
    p56_nor_69853 <= p56_nor_69853_comb;
    p56_add_69659 <= p55_add_69659;
    p56_add_69662 <= p55_add_69662;
    p56_add_69753 <= p55_add_69753;
    p56_add_69754 <= p55_add_69754;
    p56_and_69854 <= p56_and_69854_comb;
    p56_add_69875 <= p56_add_69875_comb;
    p56_add_69876 <= p56_add_69876_comb;
    p56_concat_68800 <= p55_concat_68800;
    p56_concat_69759 <= p55_concat_69759;
    p56_add_69062 <= p55_add_69062;
    p56_add_69101 <= p55_add_69101;
    p56_add_69791 <= p55_add_69791;
  end

  // ===== Pipe stage 57:
  wire [31:0] p57_add_69932_comb;
  wire [31:0] p57_and_69937_comb;
  wire [31:0] p57_add_69933_comb;
  wire [31:0] p57_add_69934_comb;
  wire [31:0] p57_add_69956_comb;
  wire [31:0] p57_nor_69936_comb;
  wire [31:0] p57_add_69958_comb;
  wire [31:0] p57_add_69959_comb;
  assign p57_add_69932_comb = (p56_add_69851 & p56_add_69726 ^ p56_nor_69853) + {p56_add_69851[5:0] ^ p56_add_69851[10:5] ^ p56_add_69851[24:19], p56_add_69851[31:27] ^ p56_add_69851[4:0] ^ p56_add_69851[18:14], p56_add_69851[26:13] ^ p56_add_69851[31:18] ^ p56_add_69851[13:0], p56_add_69851[12:6] ^ p56_add_69851[17:11] ^ p56_add_69851[31:25]};
  assign p57_and_69937_comb = p56_add_69875 & p56_add_69753;
  assign p57_add_69933_comb = p57_add_69932_comb + p56_add_69659;
  assign p57_add_69934_comb = p57_add_69933_comb + p56_add_69662;
  assign p57_add_69956_comb = (p57_and_69937_comb ^ p56_add_69875 & p56_add_69662 ^ p56_and_69854) + p56_add_69850;
  assign p57_nor_69936_comb = ~(p57_add_69934_comb | ~p56_add_69726);
  assign p57_add_69958_comb = p57_add_69956_comb + {p56_add_69875[1:0] ^ p56_add_69875[12:11] ^ p56_add_69875[21:20], p56_add_69875[31:21] ^ p56_add_69875[10:0] ^ p56_add_69875[19:9], p56_add_69875[20:12] ^ p56_add_69875[31:23] ^ p56_add_69875[8:0], p56_add_69875[11:2] ^ p56_add_69875[22:13] ^ p56_add_69875[31:22]};
  assign p57_add_69959_comb = p56_concat_68800 + p56_add_69851;

  // Registers for pipe stage 57:
  reg [31:0] p57_add_67570;
  reg [31:0] p57_add_67604;
  reg [31:0] p57_add_69851;
  reg [31:0] p57_add_69933;
  reg [31:0] p57_add_69934;
  reg [31:0] p57_nor_69936;
  reg [31:0] p57_add_69753;
  reg [31:0] p57_add_69754;
  reg [31:0] p57_add_69875;
  reg [31:0] p57_and_69937;
  reg [31:0] p57_add_69876;
  reg [31:0] p57_add_69958;
  reg [31:0] p57_add_69959;
  reg [31:0] p57_concat_69759;
  reg [31:0] p57_add_69062;
  reg [31:0] p57_add_69101;
  reg [31:0] p57_add_69791;
  always_ff @ (posedge clk) begin
    p57_add_67570 <= p56_add_67570;
    p57_add_67604 <= p56_add_67604;
    p57_add_69851 <= p56_add_69851;
    p57_add_69933 <= p57_add_69933_comb;
    p57_add_69934 <= p57_add_69934_comb;
    p57_nor_69936 <= p57_nor_69936_comb;
    p57_add_69753 <= p56_add_69753;
    p57_add_69754 <= p56_add_69754;
    p57_add_69875 <= p56_add_69875;
    p57_and_69937 <= p57_and_69937_comb;
    p57_add_69876 <= p56_add_69876;
    p57_add_69958 <= p57_add_69958_comb;
    p57_add_69959 <= p57_add_69959_comb;
    p57_concat_69759 <= p56_concat_69759;
    p57_add_69062 <= p56_add_69062;
    p57_add_69101 <= p56_add_69101;
    p57_add_69791 <= p56_add_69791;
  end

  // ===== Pipe stage 58:
  wire [31:0] p58_add_70013_comb;
  wire [31:0] p58_and_70018_comb;
  wire [31:0] p58_add_70014_comb;
  wire [31:0] p58_add_70015_comb;
  wire [31:0] p58_add_70037_comb;
  wire [31:0] p58_nor_70017_comb;
  wire [31:0] p58_add_70039_comb;
  wire [31:0] p58_add_70040_comb;
  assign p58_add_70013_comb = {p57_add_69934[5:0] ^ p57_add_69934[10:5] ^ p57_add_69934[24:19], p57_add_69934[31:27] ^ p57_add_69934[4:0] ^ p57_add_69934[18:14], p57_add_69934[26:13] ^ p57_add_69934[31:18] ^ p57_add_69934[13:0], p57_add_69934[12:6] ^ p57_add_69934[17:11] ^ p57_add_69934[31:25]} + (p57_add_69934 & p57_add_69851 ^ p57_nor_69936);
  assign p58_and_70018_comb = p57_add_69958 & p57_add_69875;
  assign p58_add_70014_comb = p58_add_70013_comb + p57_add_69754;
  assign p58_add_70015_comb = p58_add_70014_comb + p57_add_69753;
  assign p58_add_70037_comb = (p58_and_70018_comb ^ p57_add_69958 & p57_add_69753 ^ p57_and_69937) + p57_add_69933;
  assign p58_nor_70017_comb = ~(p58_add_70015_comb | ~p57_add_69851);
  assign p58_add_70039_comb = p58_add_70037_comb + {p57_add_69958[1:0] ^ p57_add_69958[12:11] ^ p57_add_69958[21:20], p57_add_69958[31:21] ^ p57_add_69958[10:0] ^ p57_add_69958[19:9], p57_add_69958[20:12] ^ p57_add_69958[31:23] ^ p57_add_69958[8:0], p57_add_69958[11:2] ^ p57_add_69958[22:13] ^ p57_add_69958[31:22]};
  assign p58_add_70040_comb = p57_concat_69759 + p57_add_69934;

  // Registers for pipe stage 58:
  reg [31:0] p58_add_67570;
  reg [31:0] p58_add_67604;
  reg [31:0] p58_add_69934;
  reg [31:0] p58_add_70014;
  reg [31:0] p58_add_70015;
  reg [31:0] p58_add_69875;
  reg [31:0] p58_nor_70017;
  reg [31:0] p58_add_69876;
  reg [31:0] p58_add_69958;
  reg [31:0] p58_and_70018;
  reg [31:0] p58_add_70039;
  reg [31:0] p58_add_69959;
  reg [31:0] p58_add_70040;
  reg [31:0] p58_add_69062;
  reg [31:0] p58_add_69101;
  reg [31:0] p58_add_69791;
  always_ff @ (posedge clk) begin
    p58_add_67570 <= p57_add_67570;
    p58_add_67604 <= p57_add_67604;
    p58_add_69934 <= p57_add_69934;
    p58_add_70014 <= p58_add_70014_comb;
    p58_add_70015 <= p58_add_70015_comb;
    p58_add_69875 <= p57_add_69875;
    p58_nor_70017 <= p58_nor_70017_comb;
    p58_add_69876 <= p57_add_69876;
    p58_add_69958 <= p57_add_69958;
    p58_and_70018 <= p58_and_70018_comb;
    p58_add_70039 <= p58_add_70039_comb;
    p58_add_69959 <= p57_add_69959;
    p58_add_70040 <= p58_add_70040_comb;
    p58_add_69062 <= p57_add_69062;
    p58_add_69101 <= p57_add_69101;
    p58_add_69791 <= p57_add_69791;
  end

  // ===== Pipe stage 59:
  wire [31:0] p59_add_70092_comb;
  wire [31:0] p59_and_70097_comb;
  wire [31:0] p59_add_70093_comb;
  wire [31:0] p59_add_70094_comb;
  wire [31:0] p59_add_70116_comb;
  wire [31:0] p59_nor_70096_comb;
  wire [31:0] p59_add_70118_comb;
  wire [31:0] p59_add_70119_comb;
  assign p59_add_70092_comb = (p58_add_70015 & p58_add_69934 ^ p58_nor_70017) + {p58_add_70015[5:0] ^ p58_add_70015[10:5] ^ p58_add_70015[24:19], p58_add_70015[31:27] ^ p58_add_70015[4:0] ^ p58_add_70015[18:14], p58_add_70015[26:13] ^ p58_add_70015[31:18] ^ p58_add_70015[13:0], p58_add_70015[12:6] ^ p58_add_70015[17:11] ^ p58_add_70015[31:25]};
  assign p59_and_70097_comb = p58_add_70039 & p58_add_69958;
  assign p59_add_70093_comb = p59_add_70092_comb + p58_add_69876;
  assign p59_add_70094_comb = p59_add_70093_comb + p58_add_69875;
  assign p59_add_70116_comb = (p59_and_70097_comb ^ p58_add_70039 & p58_add_69875 ^ p58_and_70018) + p58_add_70014;
  assign p59_nor_70096_comb = ~(p59_add_70094_comb | ~p58_add_69934);
  assign p59_add_70118_comb = p59_add_70116_comb + {p58_add_70039[1:0] ^ p58_add_70039[12:11] ^ p58_add_70039[21:20], p58_add_70039[31:21] ^ p58_add_70039[10:0] ^ p58_add_70039[19:9], p58_add_70039[20:12] ^ p58_add_70039[31:23] ^ p58_add_70039[8:0], p58_add_70039[11:2] ^ p58_add_70039[22:13] ^ p58_add_70039[31:22]};
  assign p59_add_70119_comb = p58_add_70015 + p58_add_69062;

  // Registers for pipe stage 59:
  reg [31:0] p59_add_67570;
  reg [31:0] p59_add_67604;
  reg [31:0] p59_add_70015;
  reg [31:0] p59_add_70093;
  reg [31:0] p59_add_69958;
  reg [31:0] p59_add_70094;
  reg [31:0] p59_nor_70096;
  reg [31:0] p59_add_70039;
  reg [31:0] p59_add_69959;
  reg [31:0] p59_and_70097;
  reg [31:0] p59_add_70118;
  reg [31:0] p59_add_70040;
  reg [31:0] p59_add_70119;
  reg [31:0] p59_add_69101;
  reg [31:0] p59_add_69791;
  always_ff @ (posedge clk) begin
    p59_add_67570 <= p58_add_67570;
    p59_add_67604 <= p58_add_67604;
    p59_add_70015 <= p58_add_70015;
    p59_add_70093 <= p59_add_70093_comb;
    p59_add_69958 <= p58_add_69958;
    p59_add_70094 <= p59_add_70094_comb;
    p59_nor_70096 <= p59_nor_70096_comb;
    p59_add_70039 <= p58_add_70039;
    p59_add_69959 <= p58_add_69959;
    p59_and_70097 <= p59_and_70097_comb;
    p59_add_70118 <= p59_add_70118_comb;
    p59_add_70040 <= p58_add_70040;
    p59_add_70119 <= p59_add_70119_comb;
    p59_add_69101 <= p58_add_69101;
    p59_add_69791 <= p58_add_69791;
  end

  // ===== Pipe stage 60:
  wire [31:0] p60_add_70169_comb;
  wire [31:0] p60_and_70174_comb;
  wire [31:0] p60_add_70170_comb;
  wire [31:0] p60_add_70171_comb;
  wire [31:0] p60_add_70193_comb;
  wire [31:0] p60_nor_70173_comb;
  wire [31:0] p60_add_70195_comb;
  wire [31:0] p60_add_70196_comb;
  assign p60_add_70169_comb = (p59_add_70094 & p59_add_70015 ^ p59_nor_70096) + {p59_add_70094[5:0] ^ p59_add_70094[10:5] ^ p59_add_70094[24:19], p59_add_70094[31:27] ^ p59_add_70094[4:0] ^ p59_add_70094[18:14], p59_add_70094[26:13] ^ p59_add_70094[31:18] ^ p59_add_70094[13:0], p59_add_70094[12:6] ^ p59_add_70094[17:11] ^ p59_add_70094[31:25]};
  assign p60_and_70174_comb = p59_add_70118 & p59_add_70039;
  assign p60_add_70170_comb = p60_add_70169_comb + p59_add_69959;
  assign p60_add_70171_comb = p60_add_70170_comb + p59_add_69958;
  assign p60_add_70193_comb = (p60_and_70174_comb ^ p59_add_70118 & p59_add_69958 ^ p59_and_70097) + p59_add_70093;
  assign p60_nor_70173_comb = ~(p60_add_70171_comb | ~p59_add_70015);
  assign p60_add_70195_comb = p60_add_70193_comb + {p59_add_70118[1:0] ^ p59_add_70118[12:11] ^ p59_add_70118[21:20], p59_add_70118[31:21] ^ p59_add_70118[10:0] ^ p59_add_70118[19:9], p59_add_70118[20:12] ^ p59_add_70118[31:23] ^ p59_add_70118[8:0], p59_add_70118[11:2] ^ p59_add_70118[22:13] ^ p59_add_70118[31:22]};
  assign p60_add_70196_comb = p59_add_67570 + p59_add_70094;

  // Registers for pipe stage 60:
  reg [31:0] p60_add_67604;
  reg [31:0] p60_add_70094;
  reg [31:0] p60_add_70039;
  reg [31:0] p60_add_70170;
  reg [31:0] p60_add_70171;
  reg [31:0] p60_add_70118;
  reg [31:0] p60_nor_70173;
  reg [31:0] p60_and_70174;
  reg [31:0] p60_add_70040;
  reg [31:0] p60_add_70195;
  reg [31:0] p60_add_70119;
  reg [31:0] p60_add_69101;
  reg [31:0] p60_add_70196;
  reg [31:0] p60_add_69791;
  always_ff @ (posedge clk) begin
    p60_add_67604 <= p59_add_67604;
    p60_add_70094 <= p59_add_70094;
    p60_add_70039 <= p59_add_70039;
    p60_add_70170 <= p60_add_70170_comb;
    p60_add_70171 <= p60_add_70171_comb;
    p60_add_70118 <= p59_add_70118;
    p60_nor_70173 <= p60_nor_70173_comb;
    p60_and_70174 <= p60_and_70174_comb;
    p60_add_70040 <= p59_add_70040;
    p60_add_70195 <= p60_add_70195_comb;
    p60_add_70119 <= p59_add_70119;
    p60_add_69101 <= p59_add_69101;
    p60_add_70196 <= p60_add_70196_comb;
    p60_add_69791 <= p59_add_69791;
  end

  // ===== Pipe stage 61:
  wire [31:0] p61_add_70244_comb;
  wire [31:0] p61_and_70247_comb;
  wire [31:0] p61_add_70245_comb;
  wire [31:0] p61_add_70246_comb;
  wire [31:0] p61_add_70268_comb;
  wire [31:0] p61_nor_70267_comb;
  wire [31:0] p61_add_70270_comb;
  wire [31:0] p61_add_70271_comb;
  assign p61_add_70244_comb = (p60_add_70171 & p60_add_70094 ^ p60_nor_70173) + {p60_add_70171[5:0] ^ p60_add_70171[10:5] ^ p60_add_70171[24:19], p60_add_70171[31:27] ^ p60_add_70171[4:0] ^ p60_add_70171[18:14], p60_add_70171[26:13] ^ p60_add_70171[31:18] ^ p60_add_70171[13:0], p60_add_70171[12:6] ^ p60_add_70171[17:11] ^ p60_add_70171[31:25]};
  assign p61_and_70247_comb = p60_add_70195 & p60_add_70118;
  assign p61_add_70245_comb = p61_add_70244_comb + p60_add_70040;
  assign p61_add_70246_comb = p61_add_70245_comb + p60_add_70039;
  assign p61_add_70268_comb = (p61_and_70247_comb ^ p60_add_70195 & p60_add_70039 ^ p60_and_70174) + p60_add_70170;
  assign p61_nor_70267_comb = ~(p61_add_70246_comb | ~p60_add_70094);
  assign p61_add_70270_comb = p61_add_70268_comb + {p60_add_70195[1:0] ^ p60_add_70195[12:11] ^ p60_add_70195[21:20], p60_add_70195[31:21] ^ p60_add_70195[10:0] ^ p60_add_70195[19:9], p60_add_70195[20:12] ^ p60_add_70195[31:23] ^ p60_add_70195[8:0], p60_add_70195[11:2] ^ p60_add_70195[22:13] ^ p60_add_70195[31:22]};
  assign p61_add_70271_comb = p60_add_67604 + p60_add_70171;

  // Registers for pipe stage 61:
  reg [31:0] p61_add_70171;
  reg [31:0] p61_add_70118;
  reg [31:0] p61_add_70245;
  reg [31:0] p61_add_70195;
  reg [31:0] p61_add_70246;
  reg [31:0] p61_and_70247;
  reg [31:0] p61_nor_70267;
  reg [31:0] p61_add_70270;
  reg [31:0] p61_add_70119;
  reg [31:0] p61_add_70271;
  reg [31:0] p61_add_69101;
  reg [31:0] p61_add_70196;
  reg [31:0] p61_add_69791;
  always_ff @ (posedge clk) begin
    p61_add_70171 <= p60_add_70171;
    p61_add_70118 <= p60_add_70118;
    p61_add_70245 <= p61_add_70245_comb;
    p61_add_70195 <= p60_add_70195;
    p61_add_70246 <= p61_add_70246_comb;
    p61_and_70247 <= p61_and_70247_comb;
    p61_nor_70267 <= p61_nor_70267_comb;
    p61_add_70270 <= p61_add_70270_comb;
    p61_add_70119 <= p60_add_70119;
    p61_add_70271 <= p61_add_70271_comb;
    p61_add_69101 <= p60_add_69101;
    p61_add_70196 <= p60_add_70196;
    p61_add_69791 <= p60_add_69791;
  end

  // ===== Pipe stage 62:
  wire [31:0] p62_and_70318_comb;
  wire [31:0] p62_add_70317_comb;
  wire [31:0] p62_add_70332_comb;
  wire [31:0] p62_add_70339_comb;
  wire [31:0] p62_add_70338_comb;
  wire [31:0] p62_add_70342_comb;
  wire [31:0] p62_nor_70343_comb;
  assign p62_and_70318_comb = p61_add_70270 & p61_add_70195;
  assign p62_add_70317_comb = {p61_add_70246[5:0] ^ p61_add_70246[10:5] ^ p61_add_70246[24:19], p61_add_70246[31:27] ^ p61_add_70246[4:0] ^ p61_add_70246[18:14], p61_add_70246[26:13] ^ p61_add_70246[31:18] ^ p61_add_70246[13:0], p61_add_70246[12:6] ^ p61_add_70246[17:11] ^ p61_add_70246[31:25]} + (p61_add_70246 & p61_add_70171 ^ p61_nor_70267);
  assign p62_add_70332_comb = p62_add_70317_comb + p61_add_70119;
  assign p62_add_70339_comb = (p62_and_70318_comb ^ p61_add_70270 & p61_add_70118 ^ p61_and_70247) + p61_add_70245;
  assign p62_add_70338_comb = p62_add_70332_comb + p61_add_70118;
  assign p62_add_70342_comb = p62_add_70339_comb + {p61_add_70270[1:0] ^ p61_add_70270[12:11] ^ p61_add_70270[21:20], p61_add_70270[31:21] ^ p61_add_70270[10:0] ^ p61_add_70270[19:9], p61_add_70270[20:12] ^ p61_add_70270[31:23] ^ p61_add_70270[8:0], p61_add_70270[11:2] ^ p61_add_70270[22:13] ^ p61_add_70270[31:22]};
  assign p62_nor_70343_comb = ~(p62_add_70338_comb | ~p61_add_70171);

  // Registers for pipe stage 62:
  reg [31:0] p62_add_70195;
  reg [31:0] p62_add_70246;
  reg [31:0] p62_add_70270;
  reg [31:0] p62_and_70318;
  reg [31:0] p62_add_70332;
  reg [31:0] p62_add_70338;
  reg [31:0] p62_add_70342;
  reg [31:0] p62_nor_70343;
  reg [31:0] p62_add_70271;
  reg [31:0] p62_add_69101;
  reg [31:0] p62_add_70196;
  reg [31:0] p62_add_69791;
  always_ff @ (posedge clk) begin
    p62_add_70195 <= p61_add_70195;
    p62_add_70246 <= p61_add_70246;
    p62_add_70270 <= p61_add_70270;
    p62_and_70318 <= p62_and_70318_comb;
    p62_add_70332 <= p62_add_70332_comb;
    p62_add_70338 <= p62_add_70338_comb;
    p62_add_70342 <= p62_add_70342_comb;
    p62_nor_70343 <= p62_nor_70343_comb;
    p62_add_70271 <= p61_add_70271;
    p62_add_69101 <= p61_add_69101;
    p62_add_70196 <= p61_add_70196;
    p62_add_69791 <= p61_add_69791;
  end

  // ===== Pipe stage 63:
  wire [31:0] p63_and_70385_comb;
  wire [31:0] p63_add_70406_comb;
  wire [31:0] p63_add_70407_comb;
  wire [31:0] p63_add_70409_comb;
  wire [31:0] p63_add_70410_comb;
  wire [31:0] p63_add_70411_comb;
  assign p63_and_70385_comb = p62_add_70342 & p62_add_70270;
  assign p63_add_70406_comb = {p62_add_70338[5:0] ^ p62_add_70338[10:5] ^ p62_add_70338[24:19], p62_add_70338[31:27] ^ p62_add_70338[4:0] ^ p62_add_70338[18:14], p62_add_70338[26:13] ^ p62_add_70338[31:18] ^ p62_add_70338[13:0], p62_add_70338[12:6] ^ p62_add_70338[17:11] ^ p62_add_70338[31:25]} + (p62_add_70338 & p62_add_70246 ^ p62_nor_70343);
  assign p63_add_70407_comb = (p63_and_70385_comb ^ p62_add_70342 & p62_add_70195 ^ p62_and_70318) + p62_add_70332;
  assign p63_add_70409_comb = p62_add_70196 + p63_add_70406_comb;
  assign p63_add_70410_comb = p63_add_70407_comb + {p62_add_70342[1:0] ^ p62_add_70342[12:11] ^ p62_add_70342[21:20], p62_add_70342[31:21] ^ p62_add_70342[10:0] ^ p62_add_70342[19:9], p62_add_70342[20:12] ^ p62_add_70342[31:23] ^ p62_add_70342[8:0], p62_add_70342[11:2] ^ p62_add_70342[22:13] ^ p62_add_70342[31:22]};
  assign p63_add_70411_comb = p63_add_70409_comb + p62_add_69791;

  // Registers for pipe stage 63:
  reg [31:0] p63_add_70195;
  reg [31:0] p63_add_70246;
  reg [31:0] p63_add_70270;
  reg [31:0] p63_add_70338;
  reg [31:0] p63_add_70342;
  reg [31:0] p63_and_70385;
  reg [31:0] p63_add_70410;
  reg [31:0] p63_add_70271;
  reg [31:0] p63_add_69101;
  reg [31:0] p63_add_70411;
  always_ff @ (posedge clk) begin
    p63_add_70195 <= p62_add_70195;
    p63_add_70246 <= p62_add_70246;
    p63_add_70270 <= p62_add_70270;
    p63_add_70338 <= p62_add_70338;
    p63_add_70342 <= p62_add_70342;
    p63_and_70385 <= p63_and_70385_comb;
    p63_add_70410 <= p63_add_70410_comb;
    p63_add_70271 <= p62_add_70271;
    p63_add_69101 <= p62_add_69101;
    p63_add_70411 <= p63_add_70411_comb;
  end

  // ===== Pipe stage 64:
  wire [31:0] p64_and_70432_comb;
  wire [31:0] p64_add_70446_comb;
  wire [31:0] p64_add_70465_comb;
  wire [31:0] p64_add_70473_comb;
  wire [30:0] p64_add_70487_comb;
  wire [30:0] p64_add_70489_comb;
  wire [29:0] p64_add_70491_comb;
  wire [31:0] p64_add_70476_comb;
  wire [31:0] p64_xor_70480_comb;
  wire [31:0] p64_concat_70495_comb;
  wire [31:0] p64_concat_70496_comb;
  wire [31:0] p64_concat_70497_comb;
  wire [31:0] p64_add_70498_comb;
  wire [31:0] p64_add_70499_comb;
  wire [31:0] p64_add_70479_comb;
  assign p64_and_70432_comb = p63_add_70410 & p63_add_70342;
  assign p64_add_70446_comb = p63_add_70411 + p63_add_70195;
  assign p64_add_70465_comb = (p64_and_70432_comb ^ p63_add_70410 & p63_add_70270 ^ p63_and_70385) + p63_add_70411;
  assign p64_add_70473_comb = p64_add_70465_comb + {p63_add_70410[1:0] ^ p63_add_70410[12:11] ^ p63_add_70410[21:20], p63_add_70410[31:21] ^ p63_add_70410[10:0] ^ p63_add_70410[19:9], p63_add_70410[20:12] ^ p63_add_70410[31:23] ^ p63_add_70410[8:0], p63_add_70410[11:2] ^ p63_add_70410[22:13] ^ p63_add_70410[31:22]};
  assign p64_add_70487_comb = p63_add_70410[31:1] + 31'h1e37_79b9;
  assign p64_add_70489_comb = p63_add_70342[31:1] + 31'h52a7_fa9d;
  assign p64_add_70491_comb = p64_add_70446_comb[31:2] + 30'h26c1_5a23;
  assign p64_add_70476_comb = {p64_add_70446_comb[5:0] ^ p64_add_70446_comb[10:5] ^ p64_add_70446_comb[24:19], p64_add_70446_comb[31:27] ^ p64_add_70446_comb[4:0] ^ p64_add_70446_comb[18:14], p64_add_70446_comb[26:13] ^ p64_add_70446_comb[31:18] ^ p64_add_70446_comb[13:0], p64_add_70446_comb[12:6] ^ p64_add_70446_comb[17:11] ^ p64_add_70446_comb[31:25]} + (p64_add_70446_comb & p63_add_70338 ^ ~(p64_add_70446_comb | ~p63_add_70246));
  assign p64_xor_70480_comb = p64_add_70473_comb & p63_add_70410 ^ p64_add_70473_comb & p63_add_70342 ^ p64_and_70432_comb;
  assign p64_concat_70495_comb = {p64_add_70487_comb, p63_add_70410[0]};
  assign p64_concat_70496_comb = {p64_add_70489_comb, p63_add_70342[0]};
  assign p64_concat_70497_comb = {p64_add_70491_comb, p64_add_70446_comb[1:0]};
  assign p64_add_70498_comb = p63_add_70338 + 32'h1f83_d9ab;
  assign p64_add_70499_comb = p63_add_70246 + 32'h5be0_cd19;
  assign p64_add_70479_comb = p63_add_70271 + p64_add_70476_comb;

  // Registers for pipe stage 64:
  reg [31:0] p64_add_70270;
  reg [31:0] p64_add_70473;
  reg [31:0] p64_xor_70480;
  reg [31:0] p64_concat_70495;
  reg [31:0] p64_concat_70496;
  reg [31:0] p64_concat_70497;
  reg [31:0] p64_add_70498;
  reg [31:0] p64_add_70499;
  reg [31:0] p64_add_70479;
  reg [31:0] p64_add_69101;
  always_ff @ (posedge clk) begin
    p64_add_70270 <= p63_add_70270;
    p64_add_70473 <= p64_add_70473_comb;
    p64_xor_70480 <= p64_xor_70480_comb;
    p64_concat_70495 <= p64_concat_70495_comb;
    p64_concat_70496 <= p64_concat_70496_comb;
    p64_concat_70497 <= p64_concat_70497_comb;
    p64_add_70498 <= p64_add_70498_comb;
    p64_add_70499 <= p64_add_70499_comb;
    p64_add_70479 <= p64_add_70479_comb;
    p64_add_69101 <= p63_add_69101;
  end

  // ===== Pipe stage 65:
  wire [31:0] p65_add_70537_comb;
  wire [31:0] p65_add_70540_comb;
  wire [31:0] p65_add_70541_comb;
  wire [31:0] p65_add_70543_comb;
  wire [31:0] p65_add_70544_comb;
  wire [31:0] p65_add_70545_comb;
  wire [31:0] p65_add_70546_comb;
  wire [255:0] p65_tuple_70547_comb;
  assign p65_add_70537_comb = p64_add_70479 + p64_add_69101;
  assign p65_add_70540_comb = p64_xor_70480 + {p64_add_70473[1:0] ^ p64_add_70473[12:11] ^ p64_add_70473[21:20], p64_add_70473[31:21] ^ p64_add_70473[10:0] ^ p64_add_70473[19:9], p64_add_70473[20:12] ^ p64_add_70473[31:23] ^ p64_add_70473[8:0], p64_add_70473[11:2] ^ p64_add_70473[22:13] ^ p64_add_70473[31:22]};
  assign p65_add_70541_comb = p65_add_70537_comb + 32'h6a09_e667;
  assign p65_add_70543_comb = p65_add_70537_comb + 32'h510e_527f;
  assign p65_add_70544_comb = p65_add_70540_comb + p65_add_70541_comb;
  assign p65_add_70545_comb = p64_add_70473 + 32'hbb67_ae85;
  assign p65_add_70546_comb = p65_add_70543_comb + p64_add_70270;
  assign p65_tuple_70547_comb = {p65_add_70544_comb, p65_add_70545_comb, p64_concat_70495, p64_concat_70496, p65_add_70546_comb, p64_concat_70497, p64_add_70498, p64_add_70499};

  // Registers for pipe stage 65:
  reg [255:0] p65_tuple_70547;
  always_ff @ (posedge clk) begin
    p65_tuple_70547 <= p65_tuple_70547_comb;
  end
  assign out = p65_tuple_70547;
endmodule
