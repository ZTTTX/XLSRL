module xls_test(
  input wire clk,
  input wire [511:0] message,
  output wire [255:0] out
);
  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [511:0] p0_message;
  always_ff @ (posedge clk) begin
    p0_message <= message;
  end

  // ===== Pipe stage 1:
  wire [28:0] p1_add_63010_comb;
  wire [30:0] p1_add_63014_comb;
  wire p1_bit_slice_63016_comb;
  wire [31:0] p1_concat_63033_comb;
  wire [29:0] p1_add_63040_comb;
  wire [31:0] p1_add_63047_comb;
  wire [31:0] p1_add_63048_comb;
  assign p1_add_63010_comb = p0_message[511:483] + 29'h1e6e_fdad;
  assign p1_add_63014_comb = {p1_add_63010_comb, p0_message[482:481]} + 31'h52a7_fa9d;
  assign p1_bit_slice_63016_comb = p0_message[480];
  assign p1_concat_63033_comb = {p1_add_63014_comb, p1_bit_slice_63016_comb};
  assign p1_add_63040_comb = p0_message[479:450] + 30'h242e_c78f;
  assign p1_add_63047_comb = {{p1_add_63014_comb[4:0], p1_bit_slice_63016_comb} ^ p1_add_63014_comb[9:4] ^ p1_add_63014_comb[23:18], p1_add_63014_comb[30:26] ^ {p1_add_63014_comb[3:0], p1_bit_slice_63016_comb} ^ p1_add_63014_comb[17:13], p1_add_63014_comb[25:12] ^ p1_add_63014_comb[30:17] ^ {p1_add_63014_comb[12:0], p1_bit_slice_63016_comb}, p1_add_63014_comb[11:5] ^ p1_add_63014_comb[16:10] ^ p1_add_63014_comb[30:24]} + {p1_add_63040_comb, p0_message[449:448]};
  assign p1_add_63048_comb = (p1_concat_63033_comb & 32'h510e_527f ^ ~(p1_concat_63033_comb | 32'h64fa_9773)) + p1_add_63047_comb;

  // Registers for pipe stage 1:
  reg [511:0] p1_message;
  reg [28:0] p1_add_63010;
  reg [30:0] p1_add_63014;
  reg p1_bit_slice_63016;
  reg [31:0] p1_concat_63033;
  reg [31:0] p1_add_63048;
  always_ff @ (posedge clk) begin
    p1_message <= p0_message;
    p1_add_63010 <= p1_add_63010_comb;
    p1_add_63014 <= p1_add_63014_comb;
    p1_bit_slice_63016 <= p1_bit_slice_63016_comb;
    p1_concat_63033 <= p1_concat_63033_comb;
    p1_add_63048 <= p1_add_63048_comb;
  end

  // ===== Pipe stage 2:
  wire [30:0] p2_add_63063_comb;
  wire [31:0] p2_concat_63070_comb;
  wire [31:0] p2_add_63094_comb;
  wire [31:0] p2_add_63095_comb;
  wire [31:0] p2_add_63096_comb;
  wire [31:0] p2_add_63098_comb;
  wire [29:0] p2_add_63104_comb;
  wire [31:0] p2_xor_63107_comb;
  wire [31:0] p2_concat_63110_comb;
  wire [31:0] p2_add_63127_comb;
  assign p2_add_63063_comb = p1_add_63048[31:1] + 31'h1e37_79b9;
  assign p2_concat_63070_comb = {p2_add_63063_comb, p1_add_63048[0]};
  assign p2_add_63094_comb = ({p2_add_63063_comb & p1_add_63014, p1_add_63048[0] & p1_bit_slice_63016} ^ ~(p2_concat_63070_comb | 32'haef1_ad80)) + {{p2_add_63063_comb[4:0], p1_add_63048[0]} ^ p2_add_63063_comb[9:4] ^ p2_add_63063_comb[23:18], p2_add_63063_comb[30:26] ^ {p2_add_63063_comb[3:0], p1_add_63048[0]} ^ p2_add_63063_comb[17:13], p2_add_63063_comb[25:12] ^ p2_add_63063_comb[30:17] ^ {p2_add_63063_comb[12:0], p1_add_63048[0]}, p2_add_63063_comb[11:5] ^ p2_add_63063_comb[16:10] ^ p2_add_63063_comb[30:24]};
  assign p2_add_63095_comb = p1_message[447:416] + 32'h50c6_645b;
  assign p2_add_63096_comb = p2_add_63094_comb + p2_add_63095_comb;
  assign p2_add_63098_comb = p2_add_63096_comb + 32'hbb67_ae85;
  assign p2_add_63104_comb = p1_message[415:386] + 30'h0eb1_0b89;
  assign p2_xor_63107_comb = p2_add_63098_comb & p2_concat_63070_comb ^ ~(p2_add_63098_comb | {~p1_add_63014, ~p1_bit_slice_63016});
  assign p2_concat_63110_comb = {~p2_add_63063_comb, ~p1_add_63048[0]};
  assign p2_add_63127_comb = {p1_message[390:388] ^ p1_message[401:399], p1_message[387:384] ^ p1_message[398:395] ^ p1_message[415:412], p1_message[415:405] ^ p1_message[394:384] ^ p1_message[411:401], p1_message[404:391] ^ p1_message[415:402] ^ p1_message[400:387]} + p1_message[447:416];

  // Registers for pipe stage 2:
  reg [511:0] p2_message;
  reg [28:0] p2_add_63010;
  reg [31:0] p2_concat_63033;
  reg [31:0] p2_add_63048;
  reg [31:0] p2_concat_63070;
  reg [31:0] p2_add_63098;
  reg [29:0] p2_add_63104;
  reg [31:0] p2_xor_63107;
  reg [31:0] p2_concat_63110;
  reg [31:0] p2_add_63127;
  reg [31:0] p2_add_63096;
  always_ff @ (posedge clk) begin
    p2_message <= p1_message;
    p2_add_63010 <= p1_add_63010;
    p2_concat_63033 <= p1_concat_63033;
    p2_add_63048 <= p1_add_63048;
    p2_concat_63070 <= p2_concat_63070_comb;
    p2_add_63098 <= p2_add_63098_comb;
    p2_add_63104 <= p2_add_63104_comb;
    p2_xor_63107 <= p2_xor_63107_comb;
    p2_concat_63110 <= p2_concat_63110_comb;
    p2_add_63127 <= p2_add_63127_comb;
    p2_add_63096 <= p2_add_63096_comb;
  end

  // ===== Pipe stage 3:
  wire [31:0] p3_add_63169_comb;
  wire [31:0] p3_add_63170_comb;
  wire [31:0] p3_add_63197_comb;
  wire [31:0] p3_add_63172_comb;
  wire [31:0] p3_and_63216_comb;
  wire [31:0] p3_add_63221_comb;
  wire [31:0] p3_add_63194_comb;
  wire [31:0] p3_add_63222_comb;
  assign p3_add_63169_comb = {p2_add_63098[5:0] ^ p2_add_63098[10:5] ^ p2_add_63098[24:19], p2_add_63098[31:27] ^ p2_add_63098[4:0] ^ p2_add_63098[18:14], p2_add_63098[26:13] ^ p2_add_63098[31:18] ^ p2_add_63098[13:0], p2_add_63098[12:6] ^ p2_add_63098[17:11] ^ p2_add_63098[31:25]} + {p2_add_63104, p2_message[385:384]};
  assign p3_add_63170_comb = p2_xor_63107 + p3_add_63169_comb;
  assign p3_add_63197_comb = {p2_add_63010, p2_message[482:480]} + 32'h0890_9ae5;
  assign p3_add_63172_comb = p3_add_63170_comb + 32'h6a09_e667;
  assign p3_and_63216_comb = p3_add_63197_comb & 32'h6a09_e667;
  assign p3_add_63221_comb = {p3_add_63197_comb[1:0] ^ p3_add_63197_comb[12:11] ^ p3_add_63197_comb[21:20], p3_add_63197_comb[31:21] ^ p3_add_63197_comb[10:0] ^ p3_add_63197_comb[19:9], p3_add_63197_comb[20:12] ^ p3_add_63197_comb[31:23] ^ p3_add_63197_comb[8:0], p3_add_63197_comb[11:2] ^ p3_add_63197_comb[22:13] ^ p3_add_63197_comb[31:22]} + (p3_and_63216_comb ^ p3_add_63197_comb & 32'hbb67_ae85 ^ 32'h2a01_a605);
  assign p3_add_63194_comb = {p3_add_63172_comb[5:0] ^ p3_add_63172_comb[10:5] ^ p3_add_63172_comb[24:19], p3_add_63172_comb[31:27] ^ p3_add_63172_comb[4:0] ^ p3_add_63172_comb[18:14], p3_add_63172_comb[26:13] ^ p3_add_63172_comb[31:18] ^ p3_add_63172_comb[13:0], p3_add_63172_comb[12:6] ^ p3_add_63172_comb[17:11] ^ p3_add_63172_comb[31:25]} + (p3_add_63172_comb & p2_add_63098 ^ ~(p3_add_63172_comb | p2_concat_63110));
  assign p3_add_63222_comb = p2_add_63048 + p3_add_63221_comb;

  // Registers for pipe stage 3:
  reg [511:0] p3_message;
  reg [31:0] p3_concat_63033;
  reg [31:0] p3_concat_63070;
  reg [31:0] p3_add_63098;
  reg [31:0] p3_add_63170;
  reg [31:0] p3_add_63172;
  reg [31:0] p3_add_63194;
  reg [31:0] p3_add_63197;
  reg [31:0] p3_and_63216;
  reg [31:0] p3_add_63222;
  reg [31:0] p3_add_63127;
  reg [31:0] p3_add_63096;
  always_ff @ (posedge clk) begin
    p3_message <= p2_message;
    p3_concat_63033 <= p2_concat_63033;
    p3_concat_63070 <= p2_concat_63070;
    p3_add_63098 <= p2_add_63098;
    p3_add_63170 <= p3_add_63170_comb;
    p3_add_63172 <= p3_add_63172_comb;
    p3_add_63194 <= p3_add_63194_comb;
    p3_add_63197 <= p3_add_63197_comb;
    p3_and_63216 <= p3_and_63216_comb;
    p3_add_63222 <= p3_add_63222_comb;
    p3_add_63127 <= p2_add_63127;
    p3_add_63096 <= p2_add_63096;
  end

  // ===== Pipe stage 4:
  wire [31:0] p4_and_63292_comb;
  wire [31:0] p4_add_63249_comb;
  wire [31:0] p4_add_63250_comb;
  wire [31:0] p4_add_63296_comb;
  wire [31:0] p4_add_63251_comb;
  wire [31:0] p4_add_63297_comb;
  wire [31:0] p4_add_63252_comb;
  wire [31:0] p4_and_63314_comb;
  wire [31:0] p4_add_63318_comb;
  wire [31:0] p4_add_63274_comb;
  wire [31:0] p4_add_63319_comb;
  wire [31:0] p4_add_63336_comb;
  assign p4_and_63292_comb = p3_add_63222 & p3_add_63197;
  assign p4_add_63249_comb = p3_add_63194 + 32'h3956_c25b;
  assign p4_add_63250_comb = p3_concat_63033 + p3_message[383:352];
  assign p4_add_63296_comb = {p3_add_63222[1:0] ^ p3_add_63222[12:11] ^ p3_add_63222[21:20], p3_add_63222[31:21] ^ p3_add_63222[10:0] ^ p3_add_63222[19:9], p3_add_63222[20:12] ^ p3_add_63222[31:23] ^ p3_add_63222[8:0], p3_add_63222[11:2] ^ p3_add_63222[22:13] ^ p3_add_63222[31:22]} + (p4_and_63292_comb ^ p3_add_63222 & 32'h6a09_e667 ^ p3_and_63216);
  assign p4_add_63251_comb = p4_add_63249_comb + p4_add_63250_comb;
  assign p4_add_63297_comb = p3_add_63096 + p4_add_63296_comb;
  assign p4_add_63252_comb = p3_add_63197 + p4_add_63251_comb;
  assign p4_and_63314_comb = p4_add_63297_comb & p3_add_63222;
  assign p4_add_63318_comb = {p4_add_63297_comb[1:0] ^ p4_add_63297_comb[12:11] ^ p4_add_63297_comb[21:20], p4_add_63297_comb[31:21] ^ p4_add_63297_comb[10:0] ^ p4_add_63297_comb[19:9], p4_add_63297_comb[20:12] ^ p4_add_63297_comb[31:23] ^ p4_add_63297_comb[8:0], p4_add_63297_comb[11:2] ^ p4_add_63297_comb[22:13] ^ p4_add_63297_comb[31:22]} + (p4_and_63314_comb ^ p4_add_63297_comb & p3_add_63197 ^ p4_and_63292_comb);
  assign p4_add_63274_comb = {p4_add_63252_comb[5:0] ^ p4_add_63252_comb[10:5] ^ p4_add_63252_comb[24:19], p4_add_63252_comb[31:27] ^ p4_add_63252_comb[4:0] ^ p4_add_63252_comb[18:14], p4_add_63252_comb[26:13] ^ p4_add_63252_comb[31:18] ^ p4_add_63252_comb[13:0], p4_add_63252_comb[12:6] ^ p4_add_63252_comb[17:11] ^ p4_add_63252_comb[31:25]} + (p4_add_63252_comb & p3_add_63172 ^ ~(p4_add_63252_comb | ~p3_add_63098));
  assign p4_add_63319_comb = p3_add_63170 + p4_add_63318_comb;
  assign p4_add_63336_comb = {p3_message[326:324] ^ p3_message[337:335], p3_message[323:320] ^ p3_message[334:331] ^ p3_message[351:348], p3_message[351:341] ^ p3_message[330:320] ^ p3_message[347:337], p3_message[340:327] ^ p3_message[351:338] ^ p3_message[336:323]} + p3_message[383:352];

  // Registers for pipe stage 4:
  reg [511:0] p4_message;
  reg [31:0] p4_concat_63070;
  reg [31:0] p4_add_63098;
  reg [31:0] p4_add_63172;
  reg [31:0] p4_add_63251;
  reg [31:0] p4_add_63252;
  reg [31:0] p4_add_63274;
  reg [31:0] p4_add_63222;
  reg [31:0] p4_add_63297;
  reg [31:0] p4_and_63314;
  reg [31:0] p4_add_63319;
  reg [31:0] p4_add_63336;
  reg [31:0] p4_add_63127;
  always_ff @ (posedge clk) begin
    p4_message <= p3_message;
    p4_concat_63070 <= p3_concat_63070;
    p4_add_63098 <= p3_add_63098;
    p4_add_63172 <= p3_add_63172;
    p4_add_63251 <= p4_add_63251_comb;
    p4_add_63252 <= p4_add_63252_comb;
    p4_add_63274 <= p4_add_63274_comb;
    p4_add_63222 <= p3_add_63222;
    p4_add_63297 <= p4_add_63297_comb;
    p4_and_63314 <= p4_and_63314_comb;
    p4_add_63319 <= p4_add_63319_comb;
    p4_add_63336 <= p4_add_63336_comb;
    p4_add_63127 <= p3_add_63127;
  end

  // ===== Pipe stage 5:
  wire [31:0] p5_and_63413_comb;
  wire [31:0] p5_add_63417_comb;
  wire [31:0] p5_add_63365_comb;
  wire [31:0] p5_add_63366_comb;
  wire [31:0] p5_add_63418_comb;
  wire [31:0] p5_add_63367_comb;
  wire [31:0] p5_add_63368_comb;
  wire [31:0] p5_and_63435_comb;
  wire [29:0] p5_add_63390_comb;
  wire [31:0] p5_add_63439_comb;
  wire [31:0] p5_add_63440_comb;
  wire [31:0] p5_add_63457_comb;
  wire [31:0] p5_add_63395_comb;
  wire [31:0] p5_add_63396_comb;
  assign p5_and_63413_comb = p4_add_63319 & p4_add_63297;
  assign p5_add_63417_comb = {p4_add_63319[1:0] ^ p4_add_63319[12:11] ^ p4_add_63319[21:20], p4_add_63319[31:21] ^ p4_add_63319[10:0] ^ p4_add_63319[19:9], p4_add_63319[20:12] ^ p4_add_63319[31:23] ^ p4_add_63319[8:0], p4_add_63319[11:2] ^ p4_add_63319[22:13] ^ p4_add_63319[31:22]} + (p5_and_63413_comb ^ p4_add_63319 & p4_add_63222 ^ p4_and_63314);
  assign p5_add_63365_comb = p4_add_63274 + 32'h59f1_11f1;
  assign p5_add_63366_comb = p4_concat_63070 + p4_message[351:320];
  assign p5_add_63418_comb = p4_add_63251 + p5_add_63417_comb;
  assign p5_add_63367_comb = p5_add_63365_comb + p5_add_63366_comb;
  assign p5_add_63368_comb = p4_add_63222 + p5_add_63367_comb;
  assign p5_and_63435_comb = p5_add_63418_comb & p4_add_63319;
  assign p5_add_63390_comb = p4_message[319:290] + 30'h248f_e0a9;
  assign p5_add_63439_comb = {p5_add_63418_comb[1:0] ^ p5_add_63418_comb[12:11] ^ p5_add_63418_comb[21:20], p5_add_63418_comb[31:21] ^ p5_add_63418_comb[10:0] ^ p5_add_63418_comb[19:9], p5_add_63418_comb[20:12] ^ p5_add_63418_comb[31:23] ^ p5_add_63418_comb[8:0], p5_add_63418_comb[11:2] ^ p5_add_63418_comb[22:13] ^ p5_add_63418_comb[31:22]} + (p5_and_63435_comb ^ p5_add_63418_comb & p4_add_63297 ^ p5_and_63413_comb);
  assign p5_add_63440_comb = p5_add_63367_comb + p5_add_63439_comb;
  assign p5_add_63457_comb = {p4_message[294:292] ^ p4_message[305:303], p4_message[291:288] ^ p4_message[302:299] ^ p4_message[319:316], p4_message[319:309] ^ p4_message[298:288] ^ p4_message[315:305], p4_message[308:295] ^ p4_message[319:306] ^ p4_message[304:291]} + p4_message[351:320];
  assign p5_add_63395_comb = {p5_add_63368_comb[5:0] ^ p5_add_63368_comb[10:5] ^ p5_add_63368_comb[24:19], p5_add_63368_comb[31:27] ^ p5_add_63368_comb[4:0] ^ p5_add_63368_comb[18:14], p5_add_63368_comb[26:13] ^ p5_add_63368_comb[31:18] ^ p5_add_63368_comb[13:0], p5_add_63368_comb[12:6] ^ p5_add_63368_comb[17:11] ^ p5_add_63368_comb[31:25]} + p4_add_63098;
  assign p5_add_63396_comb = (p5_add_63368_comb & p4_add_63252 ^ ~(p5_add_63368_comb | ~p4_add_63172)) + {p5_add_63390_comb, p4_message[289:288]};

  // Registers for pipe stage 5:
  reg [511:0] p5_message;
  reg [31:0] p5_add_63172;
  reg [31:0] p5_add_63252;
  reg [31:0] p5_add_63368;
  reg [31:0] p5_add_63297;
  reg [31:0] p5_add_63319;
  reg [31:0] p5_add_63418;
  reg [31:0] p5_and_63435;
  reg [31:0] p5_add_63440;
  reg [31:0] p5_add_63457;
  reg [31:0] p5_add_63336;
  reg [31:0] p5_add_63127;
  reg [31:0] p5_add_63395;
  reg [31:0] p5_add_63396;
  always_ff @ (posedge clk) begin
    p5_message <= p4_message;
    p5_add_63172 <= p4_add_63172;
    p5_add_63252 <= p4_add_63252;
    p5_add_63368 <= p5_add_63368_comb;
    p5_add_63297 <= p4_add_63297;
    p5_add_63319 <= p4_add_63319;
    p5_add_63418 <= p5_add_63418_comb;
    p5_and_63435 <= p5_and_63435_comb;
    p5_add_63440 <= p5_add_63440_comb;
    p5_add_63457 <= p5_add_63457_comb;
    p5_add_63336 <= p4_add_63336;
    p5_add_63127 <= p4_add_63127;
    p5_add_63395 <= p5_add_63395_comb;
    p5_add_63396 <= p5_add_63396_comb;
  end

  // ===== Pipe stage 6:
  wire [31:0] p6_add_63486_comb;
  wire [31:0] p6_add_63487_comb;
  wire [31:0] p6_and_63530_comb;
  wire [31:0] p6_add_63534_comb;
  wire [31:0] p6_add_63509_comb;
  wire [31:0] p6_add_63513_comb;
  wire [31:0] p6_add_63535_comb;
  wire [31:0] p6_add_63512_comb;
  wire [31:0] p6_add_63552_comb;
  assign p6_add_63486_comb = p5_add_63395 + p5_add_63396;
  assign p6_add_63487_comb = p5_add_63297 + p6_add_63486_comb;
  assign p6_and_63530_comb = p5_add_63440 & p5_add_63418;
  assign p6_add_63534_comb = {p5_add_63440[1:0] ^ p5_add_63440[12:11] ^ p5_add_63440[21:20], p5_add_63440[31:21] ^ p5_add_63440[10:0] ^ p5_add_63440[19:9], p5_add_63440[20:12] ^ p5_add_63440[31:23] ^ p5_add_63440[8:0], p5_add_63440[11:2] ^ p5_add_63440[22:13] ^ p5_add_63440[31:22]} + (p6_and_63530_comb ^ p5_add_63440 & p5_add_63319 ^ p5_and_63435);
  assign p6_add_63509_comb = {p6_add_63487_comb[5:0] ^ p6_add_63487_comb[10:5] ^ p6_add_63487_comb[24:19], p6_add_63487_comb[31:27] ^ p6_add_63487_comb[4:0] ^ p6_add_63487_comb[18:14], p6_add_63487_comb[26:13] ^ p6_add_63487_comb[31:18] ^ p6_add_63487_comb[13:0], p6_add_63487_comb[12:6] ^ p6_add_63487_comb[17:11] ^ p6_add_63487_comb[31:25]} + (p6_add_63487_comb & p5_add_63368 ^ ~(p6_add_63487_comb | ~p5_add_63252));
  assign p6_add_63513_comb = p5_add_63172 + p5_message[287:256];
  assign p6_add_63535_comb = p6_add_63486_comb + p6_add_63534_comb;
  assign p6_add_63512_comb = p6_add_63509_comb + 32'hab1c_5ed5;
  assign p6_add_63552_comb = {p5_message[230:228] ^ p5_message[241:239], p5_message[227:224] ^ p5_message[238:235] ^ p5_message[255:252], p5_message[255:245] ^ p5_message[234:224] ^ p5_message[251:241], p5_message[244:231] ^ p5_message[255:242] ^ p5_message[240:227]} + p5_message[287:256];

  // Registers for pipe stage 6:
  reg [511:0] p6_message;
  reg [31:0] p6_add_63252;
  reg [31:0] p6_add_63368;
  reg [31:0] p6_add_63487;
  reg [31:0] p6_add_63513;
  reg [31:0] p6_add_63319;
  reg [31:0] p6_add_63418;
  reg [31:0] p6_add_63440;
  reg [31:0] p6_and_63530;
  reg [31:0] p6_add_63535;
  reg [31:0] p6_add_63512;
  reg [31:0] p6_add_63552;
  reg [31:0] p6_add_63457;
  reg [31:0] p6_add_63336;
  reg [31:0] p6_add_63127;
  always_ff @ (posedge clk) begin
    p6_message <= p5_message;
    p6_add_63252 <= p5_add_63252;
    p6_add_63368 <= p5_add_63368;
    p6_add_63487 <= p6_add_63487_comb;
    p6_add_63513 <= p6_add_63513_comb;
    p6_add_63319 <= p5_add_63319;
    p6_add_63418 <= p5_add_63418;
    p6_add_63440 <= p5_add_63440;
    p6_and_63530 <= p6_and_63530_comb;
    p6_add_63535 <= p6_add_63535_comb;
    p6_add_63512 <= p6_add_63512_comb;
    p6_add_63552 <= p6_add_63552_comb;
    p6_add_63457 <= p5_add_63457;
    p6_add_63336 <= p5_add_63336;
    p6_add_63127 <= p5_add_63127;
  end

  // ===== Pipe stage 7:
  wire [31:0] p7_add_63583_comb;
  wire [31:0] p7_add_63584_comb;
  wire [31:0] p7_and_63630_comb;
  wire [28:0] p7_add_63606_comb;
  wire [31:0] p7_add_63634_comb;
  wire [31:0] p7_add_63611_comb;
  wire [31:0] p7_add_63612_comb;
  wire [31:0] p7_add_63635_comb;
  wire [31:0] p7_add_63613_comb;
  assign p7_add_63583_comb = p6_add_63512 + p6_add_63513;
  assign p7_add_63584_comb = p6_add_63319 + p7_add_63583_comb;
  assign p7_and_63630_comb = p6_add_63535 & p6_add_63440;
  assign p7_add_63606_comb = p6_message[255:227] + 29'h1b00_f553;
  assign p7_add_63634_comb = {p6_add_63535[1:0] ^ p6_add_63535[12:11] ^ p6_add_63535[21:20], p6_add_63535[31:21] ^ p6_add_63535[10:0] ^ p6_add_63535[19:9], p6_add_63535[20:12] ^ p6_add_63535[31:23] ^ p6_add_63535[8:0], p6_add_63535[11:2] ^ p6_add_63535[22:13] ^ p6_add_63535[31:22]} + (p7_and_63630_comb ^ p6_add_63535 & p6_add_63418 ^ p6_and_63530);
  assign p7_add_63611_comb = {p7_add_63584_comb[5:0] ^ p7_add_63584_comb[10:5] ^ p7_add_63584_comb[24:19], p7_add_63584_comb[31:27] ^ p7_add_63584_comb[4:0] ^ p7_add_63584_comb[18:14], p7_add_63584_comb[26:13] ^ p7_add_63584_comb[31:18] ^ p7_add_63584_comb[13:0], p7_add_63584_comb[12:6] ^ p7_add_63584_comb[17:11] ^ p7_add_63584_comb[31:25]} + p6_add_63252;
  assign p7_add_63612_comb = (p7_add_63584_comb & p6_add_63487 ^ ~(p7_add_63584_comb | ~p6_add_63368)) + {p7_add_63606_comb, p6_message[226:224]};
  assign p7_add_63635_comb = p7_add_63583_comb + p7_add_63634_comb;
  assign p7_add_63613_comb = p7_add_63611_comb + p7_add_63612_comb;

  // Registers for pipe stage 7:
  reg [511:0] p7_message;
  reg [31:0] p7_add_63368;
  reg [31:0] p7_add_63487;
  reg [31:0] p7_add_63584;
  reg [31:0] p7_add_63418;
  reg [31:0] p7_add_63440;
  reg [31:0] p7_add_63535;
  reg [31:0] p7_and_63630;
  reg [31:0] p7_add_63635;
  reg [31:0] p7_add_63552;
  reg [31:0] p7_add_63457;
  reg [31:0] p7_add_63336;
  reg [31:0] p7_add_63127;
  reg [31:0] p7_add_63613;
  always_ff @ (posedge clk) begin
    p7_message <= p6_message;
    p7_add_63368 <= p6_add_63368;
    p7_add_63487 <= p6_add_63487;
    p7_add_63584 <= p7_add_63584_comb;
    p7_add_63418 <= p6_add_63418;
    p7_add_63440 <= p6_add_63440;
    p7_add_63535 <= p6_add_63535;
    p7_and_63630 <= p7_and_63630_comb;
    p7_add_63635 <= p7_add_63635_comb;
    p7_add_63552 <= p6_add_63552;
    p7_add_63457 <= p6_add_63457;
    p7_add_63336 <= p6_add_63336;
    p7_add_63127 <= p6_add_63127;
    p7_add_63613 <= p7_add_63613_comb;
  end

  // ===== Pipe stage 8:
  wire [31:0] p8_add_63664_comb;
  wire [31:0] p8_and_63708_comb;
  wire [31:0] p8_add_63686_comb;
  wire [31:0] p8_add_63689_comb;
  wire [31:0] p8_add_63690_comb;
  wire [31:0] p8_add_63712_comb;
  wire [31:0] p8_add_63747_comb;
  wire [31:0] p8_add_63748_comb;
  wire [31:0] p8_add_63691_comb;
  wire [31:0] p8_add_63713_comb;
  wire [31:0] p8_add_63766_comb;
  wire [31:0] p8_add_63749_comb;
  assign p8_add_63664_comb = p7_add_63418 + p7_add_63613;
  assign p8_and_63708_comb = p7_add_63635 & p7_add_63535;
  assign p8_add_63686_comb = {p8_add_63664_comb[5:0] ^ p8_add_63664_comb[10:5] ^ p8_add_63664_comb[24:19], p8_add_63664_comb[31:27] ^ p8_add_63664_comb[4:0] ^ p8_add_63664_comb[18:14], p8_add_63664_comb[26:13] ^ p8_add_63664_comb[31:18] ^ p8_add_63664_comb[13:0], p8_add_63664_comb[12:6] ^ p8_add_63664_comb[17:11] ^ p8_add_63664_comb[31:25]} + (p8_add_63664_comb & p7_add_63584 ^ ~(p8_add_63664_comb | ~p7_add_63487));
  assign p8_add_63689_comb = p8_add_63686_comb + 32'h1283_5b01;
  assign p8_add_63690_comb = p7_add_63368 + p7_message[223:192];
  assign p8_add_63712_comb = {p7_add_63635[1:0] ^ p7_add_63635[12:11] ^ p7_add_63635[21:20], p7_add_63635[31:21] ^ p7_add_63635[10:0] ^ p7_add_63635[19:9], p7_add_63635[20:12] ^ p7_add_63635[31:23] ^ p7_add_63635[8:0], p7_add_63635[11:2] ^ p7_add_63635[22:13] ^ p7_add_63635[31:22]} + (p8_and_63708_comb ^ p7_add_63635 & p7_add_63440 ^ p7_and_63630);
  assign p8_add_63747_comb = {p7_message[454:452] ^ p7_message[465:463], p7_message[451:448] ^ p7_message[462:459] ^ p7_message[479:476], p7_message[479:469] ^ p7_message[458:448] ^ p7_message[475:465], p7_message[468:455] ^ p7_message[479:466] ^ p7_message[464:451]} + p7_message[511:480];
  assign p8_add_63748_comb = p7_message[223:192] + {p7_message[48:39] ^ p7_message[50:41], p7_message[38:32] ^ p7_message[40:34] ^ p7_message[63:57], p7_message[63:62] ^ p7_message[33:32] ^ p7_message[56:55], p7_message[61:49] ^ p7_message[63:51] ^ p7_message[54:42]};
  assign p8_add_63691_comb = p8_add_63689_comb + p8_add_63690_comb;
  assign p8_add_63713_comb = p7_add_63613 + p8_add_63712_comb;
  assign p8_add_63766_comb = {p7_message[166:164] ^ p7_message[177:175], p7_message[163:160] ^ p7_message[174:171] ^ p7_message[191:188], p7_message[191:181] ^ p7_message[170:160] ^ p7_message[187:177], p7_message[180:167] ^ p7_message[191:178] ^ p7_message[176:163]} + p7_message[223:192];
  assign p8_add_63749_comb = p8_add_63747_comb + p8_add_63748_comb;

  // Registers for pipe stage 8:
  reg [511:0] p8_message;
  reg [31:0] p8_add_63487;
  reg [31:0] p8_add_63584;
  reg [31:0] p8_add_63664;
  reg [31:0] p8_add_63440;
  reg [31:0] p8_add_63691;
  reg [31:0] p8_add_63535;
  reg [31:0] p8_add_63635;
  reg [31:0] p8_and_63708;
  reg [31:0] p8_add_63713;
  reg [31:0] p8_add_63766;
  reg [31:0] p8_add_63552;
  reg [31:0] p8_add_63457;
  reg [31:0] p8_add_63336;
  reg [31:0] p8_add_63127;
  reg [31:0] p8_add_63749;
  always_ff @ (posedge clk) begin
    p8_message <= p7_message;
    p8_add_63487 <= p7_add_63487;
    p8_add_63584 <= p7_add_63584;
    p8_add_63664 <= p8_add_63664_comb;
    p8_add_63440 <= p7_add_63440;
    p8_add_63691 <= p8_add_63691_comb;
    p8_add_63535 <= p7_add_63535;
    p8_add_63635 <= p7_add_63635;
    p8_and_63708 <= p8_and_63708_comb;
    p8_add_63713 <= p8_add_63713_comb;
    p8_add_63766 <= p8_add_63766_comb;
    p8_add_63552 <= p7_add_63552;
    p8_add_63457 <= p7_add_63457;
    p8_add_63336 <= p7_add_63336;
    p8_add_63127 <= p7_add_63127;
    p8_add_63749 <= p8_add_63749_comb;
  end

  // ===== Pipe stage 9:
  wire [31:0] p9_and_63855_comb;
  wire [31:0] p9_add_63799_comb;
  wire [31:0] p9_add_63862_comb;
  wire [31:0] p9_add_63944_comb;
  wire [31:0] p9_add_63925_comb;
  wire [31:0] p9_add_63926_comb;
  wire [31:0] p9_add_63863_comb;
  wire [31:0] p9_add_63945_comb;
  wire [31:0] p9_add_63927_comb;
  wire [30:0] p9_add_63821_comb;
  wire [31:0] p9_and_63880_comb;
  wire [31:0] p9_add_63826_comb;
  wire [31:0] p9_add_63827_comb;
  wire [31:0] p9_add_63828_comb;
  wire [29:0] p9_add_63834_comb;
  wire [30:0] p9_add_63857_comb;
  wire [31:0] p9_add_63885_comb;
  wire [29:0] p9_add_63889_comb;
  wire [31:0] p9_bit_slice_63884_comb;
  wire [31:0] p9_add_64000_comb;
  wire [31:0] p9_add_63980_comb;
  wire [31:0] p9_add_63981_comb;
  wire [31:0] p9_add_63829_comb;
  wire [31:0] p9_add_63831_comb;
  wire [31:0] p9_concat_63836_comb;
  wire [31:0] p9_concat_63861_comb;
  wire [31:0] p9_add_63886_comb;
  wire [31:0] p9_concat_63891_comb;
  wire [31:0] p9_bit_slice_64019_comb;
  wire [31:0] p9_add_64123_comb;
  wire [31:0] p9_add_64106_comb;
  wire [31:0] p9_add_64089_comb;
  wire [31:0] p9_add_64072_comb;
  wire [31:0] p9_add_64055_comb;
  wire [31:0] p9_add_64038_comb;
  wire [31:0] p9_add_64020_comb;
  wire [31:0] p9_add_64001_comb;
  wire [31:0] p9_add_63982_comb;
  assign p9_and_63855_comb = p8_add_63713 & p8_add_63635;
  assign p9_add_63799_comb = p8_add_63440 + p8_add_63691;
  assign p9_add_63862_comb = {p8_add_63713[1:0] ^ p8_add_63713[12:11] ^ p8_add_63713[21:20], p8_add_63713[31:21] ^ p8_add_63713[10:0] ^ p8_add_63713[19:9], p8_add_63713[20:12] ^ p8_add_63713[31:23] ^ p8_add_63713[8:0], p8_add_63713[11:2] ^ p8_add_63713[22:13] ^ p8_add_63713[31:22]} + (p9_and_63855_comb ^ p8_add_63713 & p8_add_63535 ^ p8_and_63708);
  assign p9_add_63944_comb = p8_message[159:128] + {p8_add_63749[16:7] ^ p8_add_63749[18:9], p8_add_63749[6:0] ^ p8_add_63749[8:2] ^ p8_add_63749[31:25], p8_add_63749[31:30] ^ p8_add_63749[1:0] ^ p8_add_63749[24:23], p8_add_63749[29:17] ^ p8_add_63749[31:19] ^ p8_add_63749[22:10]};
  assign p9_add_63925_comb = {p8_message[422:420] ^ p8_message[433:431], p8_message[419:416] ^ p8_message[430:427] ^ p8_message[447:444], p8_message[447:437] ^ p8_message[426:416] ^ p8_message[443:433], p8_message[436:423] ^ p8_message[447:434] ^ p8_message[432:419]} + p8_message[479:448];
  assign p9_add_63926_comb = p8_message[191:160] + {p8_message[16:7] ^ p8_message[18:9], p8_message[6:0] ^ p8_message[8:2] ^ p8_message[31:25], p8_message[31:30] ^ p8_message[1:0] ^ p8_message[24:23], p8_message[29:17] ^ p8_message[31:19] ^ p8_message[22:10]};
  assign p9_add_63863_comb = p8_add_63691 + p9_add_63862_comb;
  assign p9_add_63945_comb = p8_add_63127 + p9_add_63944_comb;
  assign p9_add_63927_comb = p9_add_63925_comb + p9_add_63926_comb;
  assign p9_add_63821_comb = p8_message[191:161] + 31'h1218_c2df;
  assign p9_and_63880_comb = p9_add_63863_comb & p8_add_63713;
  assign p9_add_63826_comb = {p9_add_63799_comb[5:0] ^ p9_add_63799_comb[10:5] ^ p9_add_63799_comb[24:19], p9_add_63799_comb[31:27] ^ p9_add_63799_comb[4:0] ^ p9_add_63799_comb[18:14], p9_add_63799_comb[26:13] ^ p9_add_63799_comb[31:18] ^ p9_add_63799_comb[13:0], p9_add_63799_comb[12:6] ^ p9_add_63799_comb[17:11] ^ p9_add_63799_comb[31:25]} + p8_add_63487;
  assign p9_add_63827_comb = (p9_add_63799_comb & p8_add_63664 ^ ~(p9_add_63799_comb | ~p8_add_63584)) + {p9_add_63821_comb, p8_message[160]};
  assign p9_add_63828_comb = p9_add_63826_comb + p9_add_63827_comb;
  assign p9_add_63834_comb = p8_message[127:98] + 30'h1caf_975d;
  assign p9_add_63857_comb = p8_message[95:65] + 31'h406f_58ff;
  assign p9_add_63885_comb = {p9_add_63863_comb[1:0] ^ p9_add_63863_comb[12:11] ^ p9_add_63863_comb[21:20], p9_add_63863_comb[31:21] ^ p9_add_63863_comb[10:0] ^ p9_add_63863_comb[19:9], p9_add_63863_comb[20:12] ^ p9_add_63863_comb[31:23] ^ p9_add_63863_comb[8:0], p9_add_63863_comb[11:2] ^ p9_add_63863_comb[22:13] ^ p9_add_63863_comb[31:22]} + (p9_and_63880_comb ^ p9_add_63863_comb & p8_add_63635 ^ p9_and_63855_comb);
  assign p9_add_63889_comb = p8_message[31:2] + 30'h3066_fc5d;
  assign p9_bit_slice_63884_comb = p8_message[63:32];
  assign p9_add_64000_comb = p8_message[95:64] + {p9_add_63945_comb[16:7] ^ p9_add_63945_comb[18:9], p9_add_63945_comb[6:0] ^ p9_add_63945_comb[8:2] ^ p9_add_63945_comb[31:25], p9_add_63945_comb[31:30] ^ p9_add_63945_comb[1:0] ^ p9_add_63945_comb[24:23], p9_add_63945_comb[29:17] ^ p9_add_63945_comb[31:19] ^ p9_add_63945_comb[22:10]};
  assign p9_add_63980_comb = {p8_message[358:356] ^ p8_message[369:367], p8_message[355:352] ^ p8_message[366:363] ^ p8_message[383:380], p8_message[383:373] ^ p8_message[362:352] ^ p8_message[379:369], p8_message[372:359] ^ p8_message[383:370] ^ p8_message[368:355]} + p8_message[415:384];
  assign p9_add_63981_comb = p8_message[127:96] + {p9_add_63927_comb[16:7] ^ p9_add_63927_comb[18:9], p9_add_63927_comb[6:0] ^ p9_add_63927_comb[8:2] ^ p9_add_63927_comb[31:25], p9_add_63927_comb[31:30] ^ p9_add_63927_comb[1:0] ^ p9_add_63927_comb[24:23], p9_add_63927_comb[29:17] ^ p9_add_63927_comb[31:19] ^ p9_add_63927_comb[22:10]};
  assign p9_add_63829_comb = p8_add_63535 + p9_add_63828_comb;
  assign p9_add_63831_comb = p8_add_63584 + p8_message[159:128];
  assign p9_concat_63836_comb = {p9_add_63834_comb, p8_message[97:96]};
  assign p9_concat_63861_comb = {p9_add_63857_comb, p8_message[64]};
  assign p9_add_63886_comb = p9_add_63828_comb + p9_add_63885_comb;
  assign p9_concat_63891_comb = {p9_add_63889_comb, p8_message[1:0]};
  assign p9_bit_slice_64019_comb = p8_message[31:0];
  assign p9_add_64123_comb = {p8_message[6:4] ^ p8_message[17:15], p8_message[3:0] ^ p8_message[14:11] ^ p8_message[31:28], p8_message[31:21] ^ p8_message[10:0] ^ p8_message[27:17], p8_message[20:7] ^ p8_message[31:18] ^ p8_message[16:3]} + p9_bit_slice_63884_comb;
  assign p9_add_64106_comb = {p8_message[38:36] ^ p8_message[49:47], p8_message[35:32] ^ p8_message[46:43] ^ p8_message[63:60], p8_message[63:53] ^ p8_message[42:32] ^ p8_message[59:49], p8_message[52:39] ^ p8_message[63:50] ^ p8_message[48:35]} + p8_message[95:64];
  assign p9_add_64089_comb = {p8_message[70:68] ^ p8_message[81:79], p8_message[67:64] ^ p8_message[78:75] ^ p8_message[95:92], p8_message[95:85] ^ p8_message[74:64] ^ p8_message[91:81], p8_message[84:71] ^ p8_message[95:82] ^ p8_message[80:67]} + p8_message[127:96];
  assign p9_add_64072_comb = {p8_message[102:100] ^ p8_message[113:111], p8_message[99:96] ^ p8_message[110:107] ^ p8_message[127:124], p8_message[127:117] ^ p8_message[106:96] ^ p8_message[123:113], p8_message[116:103] ^ p8_message[127:114] ^ p8_message[112:99]} + p8_message[159:128];
  assign p9_add_64055_comb = {p8_message[134:132] ^ p8_message[145:143], p8_message[131:128] ^ p8_message[142:139] ^ p8_message[159:156], p8_message[159:149] ^ p8_message[138:128] ^ p8_message[155:145], p8_message[148:135] ^ p8_message[159:146] ^ p8_message[144:131]} + p8_message[191:160];
  assign p9_add_64038_comb = {p8_message[198:196] ^ p8_message[209:207], p8_message[195:192] ^ p8_message[206:203] ^ p8_message[223:220], p8_message[223:213] ^ p8_message[202:192] ^ p8_message[219:209], p8_message[212:199] ^ p8_message[223:210] ^ p8_message[208:195]} + p8_message[255:224];
  assign p9_add_64020_comb = {p8_message[262:260] ^ p8_message[273:271], p8_message[259:256] ^ p8_message[270:267] ^ p8_message[287:284], p8_message[287:277] ^ p8_message[266:256] ^ p8_message[283:273], p8_message[276:263] ^ p8_message[287:274] ^ p8_message[272:259]} + p8_message[319:288];
  assign p9_add_64001_comb = p8_add_63336 + p9_add_64000_comb;
  assign p9_add_63982_comb = p9_add_63980_comb + p9_add_63981_comb;

  // Registers for pipe stage 9:
  reg [31:0] p9_add_63664;
  reg [31:0] p9_add_63799;
  reg [31:0] p9_add_63829;
  reg [31:0] p9_add_63831;
  reg [31:0] p9_add_63635;
  reg [31:0] p9_concat_63836;
  reg [31:0] p9_add_63713;
  reg [31:0] p9_concat_63861;
  reg [31:0] p9_add_63863;
  reg [31:0] p9_and_63880;
  reg [31:0] p9_bit_slice_63884;
  reg [31:0] p9_add_63886;
  reg [31:0] p9_concat_63891;
  reg [31:0] p9_bit_slice_64019;
  reg [31:0] p9_add_64123;
  reg [31:0] p9_add_64106;
  reg [31:0] p9_add_64089;
  reg [31:0] p9_add_64072;
  reg [31:0] p9_add_64055;
  reg [31:0] p9_add_63766;
  reg [31:0] p9_add_64038;
  reg [31:0] p9_add_63552;
  reg [31:0] p9_add_64020;
  reg [31:0] p9_add_63457;
  reg [31:0] p9_add_64001;
  reg [31:0] p9_add_63982;
  reg [31:0] p9_add_63945;
  reg [31:0] p9_add_63927;
  reg [31:0] p9_add_63749;
  always_ff @ (posedge clk) begin
    p9_add_63664 <= p8_add_63664;
    p9_add_63799 <= p9_add_63799_comb;
    p9_add_63829 <= p9_add_63829_comb;
    p9_add_63831 <= p9_add_63831_comb;
    p9_add_63635 <= p8_add_63635;
    p9_concat_63836 <= p9_concat_63836_comb;
    p9_add_63713 <= p8_add_63713;
    p9_concat_63861 <= p9_concat_63861_comb;
    p9_add_63863 <= p9_add_63863_comb;
    p9_and_63880 <= p9_and_63880_comb;
    p9_bit_slice_63884 <= p9_bit_slice_63884_comb;
    p9_add_63886 <= p9_add_63886_comb;
    p9_concat_63891 <= p9_concat_63891_comb;
    p9_bit_slice_64019 <= p9_bit_slice_64019_comb;
    p9_add_64123 <= p9_add_64123_comb;
    p9_add_64106 <= p9_add_64106_comb;
    p9_add_64089 <= p9_add_64089_comb;
    p9_add_64072 <= p9_add_64072_comb;
    p9_add_64055 <= p9_add_64055_comb;
    p9_add_63766 <= p8_add_63766;
    p9_add_64038 <= p9_add_64038_comb;
    p9_add_63552 <= p8_add_63552;
    p9_add_64020 <= p9_add_64020_comb;
    p9_add_63457 <= p8_add_63457;
    p9_add_64001 <= p9_add_64001_comb;
    p9_add_63982 <= p9_add_63982_comb;
    p9_add_63945 <= p9_add_63945_comb;
    p9_add_63927 <= p9_add_63927_comb;
    p9_add_63749 <= p8_add_63749;
  end

  // ===== Pipe stage 10:
  wire [31:0] p10_add_64203_comb;
  wire [31:0] p10_and_64224_comb;
  wire [31:0] p10_add_64205_comb;
  wire [31:0] p10_add_64206_comb;
  wire [31:0] p10_add_64228_comb;
  wire [31:0] p10_add_64246_comb;
  wire [31:0] p10_add_64207_comb;
  wire [31:0] p10_add_64229_comb;
  wire [31:0] p10_add_64264_comb;
  wire [31:0] p10_add_64247_comb;
  assign p10_add_64203_comb = {p9_add_63829[5:0] ^ p9_add_63829[10:5] ^ p9_add_63829[24:19], p9_add_63829[31:27] ^ p9_add_63829[4:0] ^ p9_add_63829[18:14], p9_add_63829[26:13] ^ p9_add_63829[31:18] ^ p9_add_63829[13:0], p9_add_63829[12:6] ^ p9_add_63829[17:11] ^ p9_add_63829[31:25]} + (p9_add_63829 & p9_add_63799 ^ ~(p9_add_63829 | ~p9_add_63664));
  assign p10_and_64224_comb = p9_add_63886 & p9_add_63863;
  assign p10_add_64205_comb = p10_add_64203_comb + 32'h550c_7dc3;
  assign p10_add_64206_comb = p10_add_64205_comb + p9_add_63831;
  assign p10_add_64228_comb = {p9_add_63886[1:0] ^ p9_add_63886[12:11] ^ p9_add_63886[21:20], p9_add_63886[31:21] ^ p9_add_63886[10:0] ^ p9_add_63886[19:9], p9_add_63886[20:12] ^ p9_add_63886[31:23] ^ p9_add_63886[8:0], p9_add_63886[11:2] ^ p9_add_63886[22:13] ^ p9_add_63886[31:22]} + (p10_and_64224_comb ^ p9_add_63886 & p9_add_63713 ^ p9_and_63880);
  assign p10_add_64246_comb = p9_bit_slice_64019 + {p9_add_64001[16:7] ^ p9_add_64001[18:9], p9_add_64001[6:0] ^ p9_add_64001[8:2] ^ p9_add_64001[31:25], p9_add_64001[31:30] ^ p9_add_64001[1:0] ^ p9_add_64001[24:23], p9_add_64001[29:17] ^ p9_add_64001[31:19] ^ p9_add_64001[22:10]};
  assign p10_add_64207_comb = p9_add_63635 + p10_add_64206_comb;
  assign p10_add_64229_comb = p10_add_64206_comb + p10_add_64228_comb;
  assign p10_add_64264_comb = {p9_add_63749[6:4] ^ p9_add_63749[17:15], p9_add_63749[3:0] ^ p9_add_63749[14:11] ^ p9_add_63749[31:28], p9_add_63749[31:21] ^ p9_add_63749[10:0] ^ p9_add_63749[27:17], p9_add_63749[20:7] ^ p9_add_63749[31:18] ^ p9_add_63749[16:3]} + p9_bit_slice_64019;
  assign p10_add_64247_comb = p9_add_64020 + p10_add_64246_comb;

  // Registers for pipe stage 10:
  reg [31:0] p10_add_63664;
  reg [31:0] p10_add_63799;
  reg [31:0] p10_add_63829;
  reg [31:0] p10_add_64207;
  reg [31:0] p10_concat_63836;
  reg [31:0] p10_add_63713;
  reg [31:0] p10_concat_63861;
  reg [31:0] p10_add_63863;
  reg [31:0] p10_bit_slice_63884;
  reg [31:0] p10_add_63886;
  reg [31:0] p10_and_64224;
  reg [31:0] p10_concat_63891;
  reg [31:0] p10_add_64229;
  reg [31:0] p10_add_64264;
  reg [31:0] p10_add_64123;
  reg [31:0] p10_add_64106;
  reg [31:0] p10_add_64089;
  reg [31:0] p10_add_64072;
  reg [31:0] p10_add_64055;
  reg [31:0] p10_add_63766;
  reg [31:0] p10_add_64038;
  reg [31:0] p10_add_63552;
  reg [31:0] p10_add_64247;
  reg [31:0] p10_add_63457;
  reg [31:0] p10_add_64001;
  reg [31:0] p10_add_63982;
  reg [31:0] p10_add_63945;
  reg [31:0] p10_add_63927;
  reg [31:0] p10_add_63749;
  always_ff @ (posedge clk) begin
    p10_add_63664 <= p9_add_63664;
    p10_add_63799 <= p9_add_63799;
    p10_add_63829 <= p9_add_63829;
    p10_add_64207 <= p10_add_64207_comb;
    p10_concat_63836 <= p9_concat_63836;
    p10_add_63713 <= p9_add_63713;
    p10_concat_63861 <= p9_concat_63861;
    p10_add_63863 <= p9_add_63863;
    p10_bit_slice_63884 <= p9_bit_slice_63884;
    p10_add_63886 <= p9_add_63886;
    p10_and_64224 <= p10_and_64224_comb;
    p10_concat_63891 <= p9_concat_63891;
    p10_add_64229 <= p10_add_64229_comb;
    p10_add_64264 <= p10_add_64264_comb;
    p10_add_64123 <= p9_add_64123;
    p10_add_64106 <= p9_add_64106;
    p10_add_64089 <= p9_add_64089;
    p10_add_64072 <= p9_add_64072;
    p10_add_64055 <= p9_add_64055;
    p10_add_63766 <= p9_add_63766;
    p10_add_64038 <= p9_add_64038;
    p10_add_63552 <= p9_add_63552;
    p10_add_64247 <= p10_add_64247_comb;
    p10_add_63457 <= p9_add_63457;
    p10_add_64001 <= p9_add_64001;
    p10_add_63982 <= p9_add_63982;
    p10_add_63945 <= p9_add_63945;
    p10_add_63927 <= p9_add_63927;
    p10_add_63749 <= p9_add_63749;
  end

  // ===== Pipe stage 11:
  wire [1:0] p11_bit_slice_64394_comb;
  wire [31:0] p11_add_64410_comb;
  wire [31:0] p11_add_64344_comb;
  wire [31:0] p11_add_64345_comb;
  wire [31:0] p11_add_64411_comb;
  wire [31:0] p11_add_64346_comb;
  wire [31:0] p11_add_64347_comb;
  wire [31:0] p11_and_64388_comb;
  wire [31:0] p11_add_64392_comb;
  wire [31:0] p11_add_64428_comb;
  wire [31:0] p11_add_64371_comb;
  wire [31:0] p11_add_64393_comb;
  wire [31:0] p11_add_64429_comb;
  wire [31:0] p11_add_64369_comb;
  wire [31:0] p11_add_64370_comb;
  assign p11_bit_slice_64394_comb = p10_add_63982[1:0];
  assign p11_add_64410_comb = p10_bit_slice_63884 + {p10_add_63982[16:7] ^ p10_add_63982[18:9], p10_add_63982[6:0] ^ p10_add_63982[8:2] ^ p10_add_63982[31:25], p10_add_63982[31:30] ^ p11_bit_slice_64394_comb ^ p10_add_63982[24:23], p10_add_63982[29:17] ^ p10_add_63982[31:19] ^ p10_add_63982[22:10]};
  assign p11_add_64344_comb = {p10_add_64207[5:0] ^ p10_add_64207[10:5] ^ p10_add_64207[24:19], p10_add_64207[31:27] ^ p10_add_64207[4:0] ^ p10_add_64207[18:14], p10_add_64207[26:13] ^ p10_add_64207[31:18] ^ p10_add_64207[13:0], p10_add_64207[12:6] ^ p10_add_64207[17:11] ^ p10_add_64207[31:25]} + p10_add_63664;
  assign p11_add_64345_comb = (p10_add_64207 & p10_add_63829 ^ ~(p10_add_64207 | ~p10_add_63799)) + p10_concat_63836;
  assign p11_add_64411_comb = p10_add_63457 + p11_add_64410_comb;
  assign p11_add_64346_comb = p11_add_64344_comb + p11_add_64345_comb;
  assign p11_add_64347_comb = p10_add_63713 + p11_add_64346_comb;
  assign p11_and_64388_comb = p10_add_64229 & p10_add_63886;
  assign p11_add_64392_comb = {p10_add_64229[1:0] ^ p10_add_64229[12:11] ^ p10_add_64229[21:20], p10_add_64229[31:21] ^ p10_add_64229[10:0] ^ p10_add_64229[19:9], p10_add_64229[20:12] ^ p10_add_64229[31:23] ^ p10_add_64229[8:0], p10_add_64229[11:2] ^ p10_add_64229[22:13] ^ p10_add_64229[31:22]} + (p11_and_64388_comb ^ p10_add_64229 & p10_add_63863 ^ p10_and_64224);
  assign p11_add_64428_comb = p10_add_63749 + {p11_add_64411_comb[16:7] ^ p11_add_64411_comb[18:9], p11_add_64411_comb[6:0] ^ p11_add_64411_comb[8:2] ^ p11_add_64411_comb[31:25], p11_add_64411_comb[31:30] ^ p11_add_64411_comb[1:0] ^ p11_add_64411_comb[24:23], p11_add_64411_comb[29:17] ^ p11_add_64411_comb[31:19] ^ p11_add_64411_comb[22:10]};
  assign p11_add_64371_comb = p10_add_63829 + p10_bit_slice_63884;
  assign p11_add_64393_comb = p11_add_64346_comb + p11_add_64392_comb;
  assign p11_add_64429_comb = p10_add_63552 + p11_add_64428_comb;
  assign p11_add_64369_comb = {p11_add_64347_comb[5:0] ^ p11_add_64347_comb[10:5] ^ p11_add_64347_comb[24:19], p11_add_64347_comb[31:27] ^ p11_add_64347_comb[4:0] ^ p11_add_64347_comb[18:14], p11_add_64347_comb[26:13] ^ p11_add_64347_comb[31:18] ^ p11_add_64347_comb[13:0], p11_add_64347_comb[12:6] ^ p11_add_64347_comb[17:11] ^ p11_add_64347_comb[31:25]} + p10_add_63799;
  assign p11_add_64370_comb = (p11_add_64347_comb & p10_add_64207 ^ ~(p11_add_64347_comb | ~p10_add_63829)) + p10_concat_63861;

  // Registers for pipe stage 11:
  reg [31:0] p11_add_64207;
  reg [31:0] p11_add_64347;
  reg [31:0] p11_add_63863;
  reg [31:0] p11_add_64371;
  reg [31:0] p11_add_63886;
  reg [31:0] p11_concat_63891;
  reg [31:0] p11_add_64229;
  reg [31:0] p11_and_64388;
  reg [31:0] p11_add_64393;
  reg [1:0] p11_bit_slice_64394;
  reg [31:0] p11_add_64264;
  reg [31:0] p11_add_64123;
  reg [31:0] p11_add_64106;
  reg [31:0] p11_add_64089;
  reg [31:0] p11_add_64072;
  reg [31:0] p11_add_64055;
  reg [31:0] p11_add_63766;
  reg [31:0] p11_add_64038;
  reg [31:0] p11_add_64429;
  reg [31:0] p11_add_64247;
  reg [31:0] p11_add_64411;
  reg [31:0] p11_add_64001;
  reg [31:0] p11_add_63982;
  reg [31:0] p11_add_63945;
  reg [31:0] p11_add_63927;
  reg [31:0] p11_add_63749;
  reg [31:0] p11_add_64369;
  reg [31:0] p11_add_64370;
  always_ff @ (posedge clk) begin
    p11_add_64207 <= p10_add_64207;
    p11_add_64347 <= p11_add_64347_comb;
    p11_add_63863 <= p10_add_63863;
    p11_add_64371 <= p11_add_64371_comb;
    p11_add_63886 <= p10_add_63886;
    p11_concat_63891 <= p10_concat_63891;
    p11_add_64229 <= p10_add_64229;
    p11_and_64388 <= p11_and_64388_comb;
    p11_add_64393 <= p11_add_64393_comb;
    p11_bit_slice_64394 <= p11_bit_slice_64394_comb;
    p11_add_64264 <= p10_add_64264;
    p11_add_64123 <= p10_add_64123;
    p11_add_64106 <= p10_add_64106;
    p11_add_64089 <= p10_add_64089;
    p11_add_64072 <= p10_add_64072;
    p11_add_64055 <= p10_add_64055;
    p11_add_63766 <= p10_add_63766;
    p11_add_64038 <= p10_add_64038;
    p11_add_64429 <= p11_add_64429_comb;
    p11_add_64247 <= p10_add_64247;
    p11_add_64411 <= p11_add_64411_comb;
    p11_add_64001 <= p10_add_64001;
    p11_add_63982 <= p10_add_63982;
    p11_add_63945 <= p10_add_63945;
    p11_add_63927 <= p10_add_63927;
    p11_add_63749 <= p10_add_63749;
    p11_add_64369 <= p11_add_64369_comb;
    p11_add_64370 <= p11_add_64370_comb;
  end

  // ===== Pipe stage 12:
  wire [31:0] p12_add_64486_comb;
  wire [31:0] p12_add_64550_comb;
  wire [31:0] p12_add_64487_comb;
  wire [31:0] p12_add_64551_comb;
  wire [31:0] p12_and_64528_comb;
  wire [31:0] p12_add_64532_comb;
  wire [31:0] p12_add_64509_comb;
  wire [31:0] p12_add_64568_comb;
  wire [31:0] p12_add_64533_comb;
  wire [31:0] p12_add_64511_comb;
  wire [31:0] p12_add_64569_comb;
  assign p12_add_64486_comb = p11_add_64369 + p11_add_64370;
  assign p12_add_64550_comb = p11_add_63945 + {p11_add_64429[16:7] ^ p11_add_64429[18:9], p11_add_64429[6:0] ^ p11_add_64429[8:2] ^ p11_add_64429[31:25], p11_add_64429[31:30] ^ p11_add_64429[1:0] ^ p11_add_64429[24:23], p11_add_64429[29:17] ^ p11_add_64429[31:19] ^ p11_add_64429[22:10]};
  assign p12_add_64487_comb = p11_add_63863 + p12_add_64486_comb;
  assign p12_add_64551_comb = p11_add_63766 + p12_add_64550_comb;
  assign p12_and_64528_comb = p11_add_64393 & p11_add_64229;
  assign p12_add_64532_comb = {p11_add_64393[1:0] ^ p11_add_64393[12:11] ^ p11_add_64393[21:20], p11_add_64393[31:21] ^ p11_add_64393[10:0] ^ p11_add_64393[19:9], p11_add_64393[20:12] ^ p11_add_64393[31:23] ^ p11_add_64393[8:0], p11_add_64393[11:2] ^ p11_add_64393[22:13] ^ p11_add_64393[31:22]} + (p12_and_64528_comb ^ p11_add_64393 & p11_add_63886 ^ p11_and_64388);
  assign p12_add_64509_comb = {p12_add_64487_comb[5:0] ^ p12_add_64487_comb[10:5] ^ p12_add_64487_comb[24:19], p12_add_64487_comb[31:27] ^ p12_add_64487_comb[4:0] ^ p12_add_64487_comb[18:14], p12_add_64487_comb[26:13] ^ p12_add_64487_comb[31:18] ^ p12_add_64487_comb[13:0], p12_add_64487_comb[12:6] ^ p12_add_64487_comb[17:11] ^ p12_add_64487_comb[31:25]} + (p12_add_64487_comb & p11_add_64347 ^ ~(p12_add_64487_comb | ~p11_add_64207));
  assign p12_add_64568_comb = p11_add_64001 + {p12_add_64551_comb[16:7] ^ p12_add_64551_comb[18:9], p12_add_64551_comb[6:0] ^ p12_add_64551_comb[8:2] ^ p12_add_64551_comb[31:25], p12_add_64551_comb[31:30] ^ p12_add_64551_comb[1:0] ^ p12_add_64551_comb[24:23], p12_add_64551_comb[29:17] ^ p12_add_64551_comb[31:19] ^ p12_add_64551_comb[22:10]};
  assign p12_add_64533_comb = p12_add_64486_comb + p12_add_64532_comb;
  assign p12_add_64511_comb = p12_add_64509_comb + 32'h9bdc_06a7;
  assign p12_add_64569_comb = p11_add_64072 + p12_add_64568_comb;

  // Registers for pipe stage 12:
  reg [31:0] p12_add_64207;
  reg [31:0] p12_add_64347;
  reg [31:0] p12_add_64487;
  reg [31:0] p12_add_64371;
  reg [31:0] p12_add_63886;
  reg [31:0] p12_concat_63891;
  reg [31:0] p12_add_64229;
  reg [31:0] p12_add_64393;
  reg [31:0] p12_and_64528;
  reg [31:0] p12_add_64533;
  reg [1:0] p12_bit_slice_64394;
  reg [31:0] p12_add_64511;
  reg [31:0] p12_add_64264;
  reg [31:0] p12_add_64123;
  reg [31:0] p12_add_64106;
  reg [31:0] p12_add_64089;
  reg [31:0] p12_add_64569;
  reg [31:0] p12_add_64055;
  reg [31:0] p12_add_64551;
  reg [31:0] p12_add_64038;
  reg [31:0] p12_add_64429;
  reg [31:0] p12_add_64247;
  reg [31:0] p12_add_64411;
  reg [31:0] p12_add_64001;
  reg [31:0] p12_add_63982;
  reg [31:0] p12_add_63945;
  reg [31:0] p12_add_63927;
  reg [31:0] p12_add_63749;
  always_ff @ (posedge clk) begin
    p12_add_64207 <= p11_add_64207;
    p12_add_64347 <= p11_add_64347;
    p12_add_64487 <= p12_add_64487_comb;
    p12_add_64371 <= p11_add_64371;
    p12_add_63886 <= p11_add_63886;
    p12_concat_63891 <= p11_concat_63891;
    p12_add_64229 <= p11_add_64229;
    p12_add_64393 <= p11_add_64393;
    p12_and_64528 <= p12_and_64528_comb;
    p12_add_64533 <= p12_add_64533_comb;
    p12_bit_slice_64394 <= p11_bit_slice_64394;
    p12_add_64511 <= p12_add_64511_comb;
    p12_add_64264 <= p11_add_64264;
    p12_add_64123 <= p11_add_64123;
    p12_add_64106 <= p11_add_64106;
    p12_add_64089 <= p11_add_64089;
    p12_add_64569 <= p12_add_64569_comb;
    p12_add_64055 <= p11_add_64055;
    p12_add_64551 <= p12_add_64551_comb;
    p12_add_64038 <= p11_add_64038;
    p12_add_64429 <= p11_add_64429;
    p12_add_64247 <= p11_add_64247;
    p12_add_64411 <= p11_add_64411;
    p12_add_64001 <= p11_add_64001;
    p12_add_63982 <= p11_add_63982;
    p12_add_63945 <= p11_add_63945;
    p12_add_63927 <= p11_add_63927;
    p12_add_63749 <= p11_add_63749;
  end

  // ===== Pipe stage 13:
  wire [31:0] p13_add_64626_comb;
  wire [31:0] p13_add_64627_comb;
  wire [31:0] p13_and_64669_comb;
  wire [31:0] p13_add_64673_comb;
  wire [31:0] p13_add_64691_comb;
  wire [31:0] p13_add_64649_comb;
  wire [31:0] p13_add_64650_comb;
  wire [31:0] p13_add_64652_comb;
  wire [31:0] p13_add_64674_comb;
  wire [31:0] p13_add_64709_comb;
  wire [31:0] p13_add_64692_comb;
  wire [31:0] p13_add_64651_comb;
  assign p13_add_64626_comb = p12_add_64511 + p12_add_64371;
  assign p13_add_64627_comb = p12_add_63886 + p13_add_64626_comb;
  assign p13_and_64669_comb = p12_add_64533 & p12_add_64393;
  assign p13_add_64673_comb = {p12_add_64533[1:0] ^ p12_add_64533[12:11] ^ p12_add_64533[21:20], p12_add_64533[31:21] ^ p12_add_64533[10:0] ^ p12_add_64533[19:9], p12_add_64533[20:12] ^ p12_add_64533[31:23] ^ p12_add_64533[8:0], p12_add_64533[11:2] ^ p12_add_64533[22:13] ^ p12_add_64533[31:22]} + (p13_and_64669_comb ^ p12_add_64533 & p12_add_64229 ^ p12_and_64528);
  assign p13_add_64691_comb = p12_add_64247 + {p12_add_64569[16:7] ^ p12_add_64569[18:9], p12_add_64569[6:0] ^ p12_add_64569[8:2] ^ p12_add_64569[31:25], p12_add_64569[31:30] ^ p12_add_64569[1:0] ^ p12_add_64569[24:23], p12_add_64569[29:17] ^ p12_add_64569[31:19] ^ p12_add_64569[22:10]};
  assign p13_add_64649_comb = {p13_add_64627_comb[5:0] ^ p13_add_64627_comb[10:5] ^ p13_add_64627_comb[24:19], p13_add_64627_comb[31:27] ^ p13_add_64627_comb[4:0] ^ p13_add_64627_comb[18:14], p13_add_64627_comb[26:13] ^ p13_add_64627_comb[31:18] ^ p13_add_64627_comb[13:0], p13_add_64627_comb[12:6] ^ p13_add_64627_comb[17:11] ^ p13_add_64627_comb[31:25]} + p12_add_64207;
  assign p13_add_64650_comb = (p13_add_64627_comb & p12_add_64487 ^ ~(p13_add_64627_comb | ~p12_add_64347)) + p12_concat_63891;
  assign p13_add_64652_comb = p12_add_64347 + p12_add_63749;
  assign p13_add_64674_comb = p13_add_64626_comb + p13_add_64673_comb;
  assign p13_add_64709_comb = {p12_add_63927[6:4] ^ p12_add_63927[17:15], p12_add_63927[3:0] ^ p12_add_63927[14:11] ^ p12_add_63927[31:28], p12_add_63927[31:21] ^ p12_add_63927[10:0] ^ p12_add_63927[27:17], p12_add_63927[20:7] ^ p12_add_63927[31:18] ^ p12_add_63927[16:3]} + p12_add_63749;
  assign p13_add_64692_comb = p12_add_64106 + p13_add_64691_comb;
  assign p13_add_64651_comb = p13_add_64649_comb + p13_add_64650_comb;

  // Registers for pipe stage 13:
  reg [31:0] p13_add_64487;
  reg [31:0] p13_add_64627;
  reg [31:0] p13_add_64229;
  reg [31:0] p13_add_64652;
  reg [31:0] p13_add_64393;
  reg [31:0] p13_add_64533;
  reg [31:0] p13_and_64669;
  reg [31:0] p13_add_64674;
  reg [1:0] p13_bit_slice_64394;
  reg [31:0] p13_add_64709;
  reg [31:0] p13_add_64264;
  reg [31:0] p13_add_64123;
  reg [31:0] p13_add_64692;
  reg [31:0] p13_add_64089;
  reg [31:0] p13_add_64569;
  reg [31:0] p13_add_64055;
  reg [31:0] p13_add_64551;
  reg [31:0] p13_add_64038;
  reg [31:0] p13_add_64429;
  reg [31:0] p13_add_64247;
  reg [31:0] p13_add_64411;
  reg [31:0] p13_add_64001;
  reg [31:0] p13_add_63982;
  reg [31:0] p13_add_63945;
  reg [31:0] p13_add_63927;
  reg [31:0] p13_add_64651;
  always_ff @ (posedge clk) begin
    p13_add_64487 <= p12_add_64487;
    p13_add_64627 <= p13_add_64627_comb;
    p13_add_64229 <= p12_add_64229;
    p13_add_64652 <= p13_add_64652_comb;
    p13_add_64393 <= p12_add_64393;
    p13_add_64533 <= p12_add_64533;
    p13_and_64669 <= p13_and_64669_comb;
    p13_add_64674 <= p13_add_64674_comb;
    p13_bit_slice_64394 <= p12_bit_slice_64394;
    p13_add_64709 <= p13_add_64709_comb;
    p13_add_64264 <= p12_add_64264;
    p13_add_64123 <= p12_add_64123;
    p13_add_64692 <= p13_add_64692_comb;
    p13_add_64089 <= p12_add_64089;
    p13_add_64569 <= p12_add_64569;
    p13_add_64055 <= p12_add_64055;
    p13_add_64551 <= p12_add_64551;
    p13_add_64038 <= p12_add_64038;
    p13_add_64429 <= p12_add_64429;
    p13_add_64247 <= p12_add_64247;
    p13_add_64411 <= p12_add_64411;
    p13_add_64001 <= p12_add_64001;
    p13_add_63982 <= p12_add_63982;
    p13_add_63945 <= p12_add_63945;
    p13_add_63927 <= p12_add_63927;
    p13_add_64651 <= p13_add_64651_comb;
  end

  // ===== Pipe stage 14:
  wire [31:0] p14_add_64762_comb;
  wire [31:0] p14_and_64804_comb;
  wire [31:0] p14_add_64784_comb;
  wire [31:0] p14_add_64786_comb;
  wire [31:0] p14_add_64808_comb;
  wire [31:0] p14_add_64787_comb;
  wire [31:0] p14_add_64809_comb;
  assign p14_add_64762_comb = p13_add_64229 + p13_add_64651;
  assign p14_and_64804_comb = p13_add_64674 & p13_add_64533;
  assign p14_add_64784_comb = {p14_add_64762_comb[5:0] ^ p14_add_64762_comb[10:5] ^ p14_add_64762_comb[24:19], p14_add_64762_comb[31:27] ^ p14_add_64762_comb[4:0] ^ p14_add_64762_comb[18:14], p14_add_64762_comb[26:13] ^ p14_add_64762_comb[31:18] ^ p14_add_64762_comb[13:0], p14_add_64762_comb[12:6] ^ p14_add_64762_comb[17:11] ^ p14_add_64762_comb[31:25]} + (p14_add_64762_comb & p13_add_64627 ^ ~(p14_add_64762_comb | ~p13_add_64487));
  assign p14_add_64786_comb = p14_add_64784_comb + 32'he49b_69c1;
  assign p14_add_64808_comb = {p13_add_64674[1:0] ^ p13_add_64674[12:11] ^ p13_add_64674[21:20], p13_add_64674[31:21] ^ p13_add_64674[10:0] ^ p13_add_64674[19:9], p13_add_64674[20:12] ^ p13_add_64674[31:23] ^ p13_add_64674[8:0], p13_add_64674[11:2] ^ p13_add_64674[22:13] ^ p13_add_64674[31:22]} + (p14_and_64804_comb ^ p13_add_64674 & p13_add_64393 ^ p13_and_64669);
  assign p14_add_64787_comb = p14_add_64786_comb + p13_add_64652;
  assign p14_add_64809_comb = p13_add_64651 + p14_add_64808_comb;

  // Registers for pipe stage 14:
  reg [31:0] p14_add_64487;
  reg [31:0] p14_add_64627;
  reg [31:0] p14_add_64762;
  reg [31:0] p14_add_64393;
  reg [31:0] p14_add_64787;
  reg [31:0] p14_add_64533;
  reg [31:0] p14_add_64674;
  reg [1:0] p14_bit_slice_64394;
  reg [31:0] p14_and_64804;
  reg [31:0] p14_add_64809;
  reg [31:0] p14_add_64709;
  reg [31:0] p14_add_64264;
  reg [31:0] p14_add_64123;
  reg [31:0] p14_add_64692;
  reg [31:0] p14_add_64089;
  reg [31:0] p14_add_64569;
  reg [31:0] p14_add_64055;
  reg [31:0] p14_add_64551;
  reg [31:0] p14_add_64038;
  reg [31:0] p14_add_64429;
  reg [31:0] p14_add_64247;
  reg [31:0] p14_add_64411;
  reg [31:0] p14_add_64001;
  reg [31:0] p14_add_63982;
  reg [31:0] p14_add_63945;
  reg [31:0] p14_add_63927;
  always_ff @ (posedge clk) begin
    p14_add_64487 <= p13_add_64487;
    p14_add_64627 <= p13_add_64627;
    p14_add_64762 <= p14_add_64762_comb;
    p14_add_64393 <= p13_add_64393;
    p14_add_64787 <= p14_add_64787_comb;
    p14_add_64533 <= p13_add_64533;
    p14_add_64674 <= p13_add_64674;
    p14_bit_slice_64394 <= p13_bit_slice_64394;
    p14_and_64804 <= p14_and_64804_comb;
    p14_add_64809 <= p14_add_64809_comb;
    p14_add_64709 <= p13_add_64709;
    p14_add_64264 <= p13_add_64264;
    p14_add_64123 <= p13_add_64123;
    p14_add_64692 <= p13_add_64692;
    p14_add_64089 <= p13_add_64089;
    p14_add_64569 <= p13_add_64569;
    p14_add_64055 <= p13_add_64055;
    p14_add_64551 <= p13_add_64551;
    p14_add_64038 <= p13_add_64038;
    p14_add_64429 <= p13_add_64429;
    p14_add_64247 <= p13_add_64247;
    p14_add_64411 <= p13_add_64411;
    p14_add_64001 <= p13_add_64001;
    p14_add_63982 <= p13_add_63982;
    p14_add_63945 <= p13_add_63945;
    p14_add_63927 <= p13_add_63927;
  end

  // ===== Pipe stage 15:
  wire [31:0] p15_and_64912_comb;
  wire [31:0] p15_add_64862_comb;
  wire [31:0] p15_add_64916_comb;
  wire [31:0] p15_add_64917_comb;
  wire [30:0] p15_add_64884_comb;
  wire [31:0] p15_and_64934_comb;
  wire [31:0] p15_add_64889_comb;
  wire [31:0] p15_add_64890_comb;
  wire [31:0] p15_add_64891_comb;
  wire [31:0] p15_add_64938_comb;
  wire [31:0] p15_add_64892_comb;
  wire [30:0] p15_add_64895_comb;
  wire [31:0] p15_add_64939_comb;
  assign p15_and_64912_comb = p14_add_64809 & p14_add_64674;
  assign p15_add_64862_comb = p14_add_64393 + p14_add_64787;
  assign p15_add_64916_comb = {p14_add_64809[1:0] ^ p14_add_64809[12:11] ^ p14_add_64809[21:20], p14_add_64809[31:21] ^ p14_add_64809[10:0] ^ p14_add_64809[19:9], p14_add_64809[20:12] ^ p14_add_64809[31:23] ^ p14_add_64809[8:0], p14_add_64809[11:2] ^ p14_add_64809[22:13] ^ p14_add_64809[31:22]} + (p15_and_64912_comb ^ p14_add_64809 & p14_add_64533 ^ p14_and_64804);
  assign p15_add_64917_comb = p14_add_64787 + p15_add_64916_comb;
  assign p15_add_64884_comb = p14_add_63927[31:1] + 31'h77df_23c3;
  assign p15_and_64934_comb = p15_add_64917_comb & p14_add_64809;
  assign p15_add_64889_comb = {p15_add_64862_comb[5:0] ^ p15_add_64862_comb[10:5] ^ p15_add_64862_comb[24:19], p15_add_64862_comb[31:27] ^ p15_add_64862_comb[4:0] ^ p15_add_64862_comb[18:14], p15_add_64862_comb[26:13] ^ p15_add_64862_comb[31:18] ^ p15_add_64862_comb[13:0], p15_add_64862_comb[12:6] ^ p15_add_64862_comb[17:11] ^ p15_add_64862_comb[31:25]} + p14_add_64487;
  assign p15_add_64890_comb = (p15_add_64862_comb & p14_add_64762 ^ ~(p15_add_64862_comb | ~p14_add_64627)) + {p15_add_64884_comb, p14_add_63927[0]};
  assign p15_add_64891_comb = p15_add_64889_comb + p15_add_64890_comb;
  assign p15_add_64938_comb = {p15_add_64917_comb[1:0] ^ p15_add_64917_comb[12:11] ^ p15_add_64917_comb[21:20], p15_add_64917_comb[31:21] ^ p15_add_64917_comb[10:0] ^ p15_add_64917_comb[19:9], p15_add_64917_comb[20:12] ^ p15_add_64917_comb[31:23] ^ p15_add_64917_comb[8:0], p15_add_64917_comb[11:2] ^ p15_add_64917_comb[22:13] ^ p15_add_64917_comb[31:22]} + (p15_and_64934_comb ^ p15_add_64917_comb & p14_add_64674 ^ p15_and_64912_comb);
  assign p15_add_64892_comb = p14_add_64533 + p15_add_64891_comb;
  assign p15_add_64895_comb = p14_add_63945[31:1] + 31'h07e0_cee3;
  assign p15_add_64939_comb = p15_add_64891_comb + p15_add_64938_comb;

  // Registers for pipe stage 15:
  reg [31:0] p15_add_64627;
  reg [31:0] p15_add_64762;
  reg [31:0] p15_add_64862;
  reg [31:0] p15_add_64892;
  reg [30:0] p15_add_64895;
  reg [31:0] p15_add_64674;
  reg [1:0] p15_bit_slice_64394;
  reg [31:0] p15_add_64809;
  reg [31:0] p15_add_64917;
  reg [31:0] p15_and_64934;
  reg [31:0] p15_add_64939;
  reg [31:0] p15_add_64709;
  reg [31:0] p15_add_64264;
  reg [31:0] p15_add_64123;
  reg [31:0] p15_add_64692;
  reg [31:0] p15_add_64089;
  reg [31:0] p15_add_64569;
  reg [31:0] p15_add_64055;
  reg [31:0] p15_add_64551;
  reg [31:0] p15_add_64038;
  reg [31:0] p15_add_64429;
  reg [31:0] p15_add_64247;
  reg [31:0] p15_add_64411;
  reg [31:0] p15_add_64001;
  reg [31:0] p15_add_63982;
  reg [31:0] p15_add_63945;
  reg [31:0] p15_add_63927;
  always_ff @ (posedge clk) begin
    p15_add_64627 <= p14_add_64627;
    p15_add_64762 <= p14_add_64762;
    p15_add_64862 <= p15_add_64862_comb;
    p15_add_64892 <= p15_add_64892_comb;
    p15_add_64895 <= p15_add_64895_comb;
    p15_add_64674 <= p14_add_64674;
    p15_bit_slice_64394 <= p14_bit_slice_64394;
    p15_add_64809 <= p14_add_64809;
    p15_add_64917 <= p15_add_64917_comb;
    p15_and_64934 <= p15_and_64934_comb;
    p15_add_64939 <= p15_add_64939_comb;
    p15_add_64709 <= p14_add_64709;
    p15_add_64264 <= p14_add_64264;
    p15_add_64123 <= p14_add_64123;
    p15_add_64692 <= p14_add_64692;
    p15_add_64089 <= p14_add_64089;
    p15_add_64569 <= p14_add_64569;
    p15_add_64055 <= p14_add_64055;
    p15_add_64551 <= p14_add_64551;
    p15_add_64038 <= p14_add_64038;
    p15_add_64429 <= p14_add_64429;
    p15_add_64247 <= p14_add_64247;
    p15_add_64411 <= p14_add_64411;
    p15_add_64001 <= p14_add_64001;
    p15_add_63982 <= p14_add_63982;
    p15_add_63945 <= p14_add_63945;
    p15_add_63927 <= p14_add_63927;
  end

  // ===== Pipe stage 16:
  wire [31:0] p16_add_65017_comb;
  wire [31:0] p16_add_65018_comb;
  wire [31:0] p16_add_65019_comb;
  wire [31:0] p16_add_65020_comb;
  wire [31:0] p16_and_65065_comb;
  wire [29:0] p16_add_65042_comb;
  wire [31:0] p16_add_65069_comb;
  wire [31:0] p16_add_65048_comb;
  wire [31:0] p16_add_65070_comb;
  wire [31:0] p16_add_65046_comb;
  wire [31:0] p16_add_65047_comb;
  assign p16_add_65017_comb = {p15_add_64892[5:0] ^ p15_add_64892[10:5] ^ p15_add_64892[24:19], p15_add_64892[31:27] ^ p15_add_64892[4:0] ^ p15_add_64892[18:14], p15_add_64892[26:13] ^ p15_add_64892[31:18] ^ p15_add_64892[13:0], p15_add_64892[12:6] ^ p15_add_64892[17:11] ^ p15_add_64892[31:25]} + p15_add_64627;
  assign p16_add_65018_comb = (p15_add_64892 & p15_add_64862 ^ ~(p15_add_64892 | ~p15_add_64762)) + {p15_add_64895, p15_add_63945[0]};
  assign p16_add_65019_comb = p16_add_65017_comb + p16_add_65018_comb;
  assign p16_add_65020_comb = p15_add_64674 + p16_add_65019_comb;
  assign p16_and_65065_comb = p15_add_64939 & p15_add_64917;
  assign p16_add_65042_comb = p15_add_63982[31:2] + 30'h0903_2873;
  assign p16_add_65069_comb = {p15_add_64939[1:0] ^ p15_add_64939[12:11] ^ p15_add_64939[21:20], p15_add_64939[31:21] ^ p15_add_64939[10:0] ^ p15_add_64939[19:9], p15_add_64939[20:12] ^ p15_add_64939[31:23] ^ p15_add_64939[8:0], p15_add_64939[11:2] ^ p15_add_64939[22:13] ^ p15_add_64939[31:22]} + (p16_and_65065_comb ^ p15_add_64939 & p15_add_64809 ^ p15_and_64934);
  assign p16_add_65048_comb = p15_add_64862 + p15_add_64001;
  assign p16_add_65070_comb = p16_add_65019_comb + p16_add_65069_comb;
  assign p16_add_65046_comb = {p16_add_65020_comb[5:0] ^ p16_add_65020_comb[10:5] ^ p16_add_65020_comb[24:19], p16_add_65020_comb[31:27] ^ p16_add_65020_comb[4:0] ^ p16_add_65020_comb[18:14], p16_add_65020_comb[26:13] ^ p16_add_65020_comb[31:18] ^ p16_add_65020_comb[13:0], p16_add_65020_comb[12:6] ^ p16_add_65020_comb[17:11] ^ p16_add_65020_comb[31:25]} + p15_add_64762;
  assign p16_add_65047_comb = (p16_add_65020_comb & p15_add_64892 ^ ~(p16_add_65020_comb | ~p15_add_64862)) + {p16_add_65042_comb, p15_bit_slice_64394};

  // Registers for pipe stage 16:
  reg [31:0] p16_add_64892;
  reg [31:0] p16_add_65020;
  reg [31:0] p16_add_64809;
  reg [31:0] p16_add_65048;
  reg [31:0] p16_add_64917;
  reg [31:0] p16_add_64939;
  reg [31:0] p16_and_65065;
  reg [31:0] p16_add_65070;
  reg [31:0] p16_add_64709;
  reg [31:0] p16_add_64264;
  reg [31:0] p16_add_64123;
  reg [31:0] p16_add_64692;
  reg [31:0] p16_add_64089;
  reg [31:0] p16_add_64569;
  reg [31:0] p16_add_64055;
  reg [31:0] p16_add_64551;
  reg [31:0] p16_add_64038;
  reg [31:0] p16_add_64429;
  reg [31:0] p16_add_64247;
  reg [31:0] p16_add_64411;
  reg [31:0] p16_add_64001;
  reg [31:0] p16_add_65046;
  reg [31:0] p16_add_65047;
  reg [31:0] p16_add_63982;
  reg [31:0] p16_add_63945;
  reg [31:0] p16_add_63927;
  always_ff @ (posedge clk) begin
    p16_add_64892 <= p15_add_64892;
    p16_add_65020 <= p16_add_65020_comb;
    p16_add_64809 <= p15_add_64809;
    p16_add_65048 <= p16_add_65048_comb;
    p16_add_64917 <= p15_add_64917;
    p16_add_64939 <= p15_add_64939;
    p16_and_65065 <= p16_and_65065_comb;
    p16_add_65070 <= p16_add_65070_comb;
    p16_add_64709 <= p15_add_64709;
    p16_add_64264 <= p15_add_64264;
    p16_add_64123 <= p15_add_64123;
    p16_add_64692 <= p15_add_64692;
    p16_add_64089 <= p15_add_64089;
    p16_add_64569 <= p15_add_64569;
    p16_add_64055 <= p15_add_64055;
    p16_add_64551 <= p15_add_64551;
    p16_add_64038 <= p15_add_64038;
    p16_add_64429 <= p15_add_64429;
    p16_add_64247 <= p15_add_64247;
    p16_add_64411 <= p15_add_64411;
    p16_add_64001 <= p15_add_64001;
    p16_add_65046 <= p16_add_65046_comb;
    p16_add_65047 <= p16_add_65047_comb;
    p16_add_63982 <= p15_add_63982;
    p16_add_63945 <= p15_add_63945;
    p16_add_63927 <= p15_add_63927;
  end

  // ===== Pipe stage 17:
  wire [31:0] p17_add_65123_comb;
  wire [31:0] p17_add_65124_comb;
  wire [31:0] p17_and_65165_comb;
  wire [31:0] p17_add_65169_comb;
  wire [31:0] p17_add_65146_comb;
  wire [31:0] p17_add_65170_comb;
  wire [31:0] p17_add_65148_comb;
  assign p17_add_65123_comb = p16_add_65046 + p16_add_65047;
  assign p17_add_65124_comb = p16_add_64809 + p17_add_65123_comb;
  assign p17_and_65165_comb = p16_add_65070 & p16_add_64939;
  assign p17_add_65169_comb = {p16_add_65070[1:0] ^ p16_add_65070[12:11] ^ p16_add_65070[21:20], p16_add_65070[31:21] ^ p16_add_65070[10:0] ^ p16_add_65070[19:9], p16_add_65070[20:12] ^ p16_add_65070[31:23] ^ p16_add_65070[8:0], p16_add_65070[11:2] ^ p16_add_65070[22:13] ^ p16_add_65070[31:22]} + (p17_and_65165_comb ^ p16_add_65070 & p16_add_64917 ^ p16_and_65065);
  assign p17_add_65146_comb = {p17_add_65124_comb[5:0] ^ p17_add_65124_comb[10:5] ^ p17_add_65124_comb[24:19], p17_add_65124_comb[31:27] ^ p17_add_65124_comb[4:0] ^ p17_add_65124_comb[18:14], p17_add_65124_comb[26:13] ^ p17_add_65124_comb[31:18] ^ p17_add_65124_comb[13:0], p17_add_65124_comb[12:6] ^ p17_add_65124_comb[17:11] ^ p17_add_65124_comb[31:25]} + (p17_add_65124_comb & p16_add_65020 ^ ~(p17_add_65124_comb | ~p16_add_64892));
  assign p17_add_65170_comb = p17_add_65123_comb + p17_add_65169_comb;
  assign p17_add_65148_comb = p17_add_65146_comb + 32'h2de9_2c6f;

  // Registers for pipe stage 17:
  reg [31:0] p17_add_64892;
  reg [31:0] p17_add_65020;
  reg [31:0] p17_add_65124;
  reg [31:0] p17_add_65048;
  reg [31:0] p17_add_64917;
  reg [31:0] p17_add_64939;
  reg [31:0] p17_add_65070;
  reg [31:0] p17_and_65165;
  reg [31:0] p17_add_65170;
  reg [31:0] p17_add_65148;
  reg [31:0] p17_add_64709;
  reg [31:0] p17_add_64264;
  reg [31:0] p17_add_64123;
  reg [31:0] p17_add_64692;
  reg [31:0] p17_add_64089;
  reg [31:0] p17_add_64569;
  reg [31:0] p17_add_64055;
  reg [31:0] p17_add_64551;
  reg [31:0] p17_add_64038;
  reg [31:0] p17_add_64429;
  reg [31:0] p17_add_64247;
  reg [31:0] p17_add_64411;
  reg [31:0] p17_add_64001;
  reg [31:0] p17_add_63982;
  reg [31:0] p17_add_63945;
  reg [31:0] p17_add_63927;
  always_ff @ (posedge clk) begin
    p17_add_64892 <= p16_add_64892;
    p17_add_65020 <= p16_add_65020;
    p17_add_65124 <= p17_add_65124_comb;
    p17_add_65048 <= p16_add_65048;
    p17_add_64917 <= p16_add_64917;
    p17_add_64939 <= p16_add_64939;
    p17_add_65070 <= p16_add_65070;
    p17_and_65165 <= p17_and_65165_comb;
    p17_add_65170 <= p17_add_65170_comb;
    p17_add_65148 <= p17_add_65148_comb;
    p17_add_64709 <= p16_add_64709;
    p17_add_64264 <= p16_add_64264;
    p17_add_64123 <= p16_add_64123;
    p17_add_64692 <= p16_add_64692;
    p17_add_64089 <= p16_add_64089;
    p17_add_64569 <= p16_add_64569;
    p17_add_64055 <= p16_add_64055;
    p17_add_64551 <= p16_add_64551;
    p17_add_64038 <= p16_add_64038;
    p17_add_64429 <= p16_add_64429;
    p17_add_64247 <= p16_add_64247;
    p17_add_64411 <= p16_add_64411;
    p17_add_64001 <= p16_add_64001;
    p17_add_63982 <= p16_add_63982;
    p17_add_63945 <= p16_add_63945;
    p17_add_63927 <= p16_add_63927;
  end

  // ===== Pipe stage 18:
  wire [31:0] p18_add_65223_comb;
  wire [31:0] p18_add_65224_comb;
  wire [31:0] p18_and_65270_comb;
  wire [30:0] p18_add_65246_comb;
  wire [31:0] p18_add_65274_comb;
  wire [31:0] p18_add_65251_comb;
  wire [31:0] p18_add_65252_comb;
  wire [31:0] p18_add_65275_comb;
  wire [31:0] p18_add_65253_comb;
  assign p18_add_65223_comb = p17_add_65148 + p17_add_65048;
  assign p18_add_65224_comb = p17_add_64917 + p18_add_65223_comb;
  assign p18_and_65270_comb = p17_add_65170 & p17_add_65070;
  assign p18_add_65246_comb = p17_add_64411[31:1] + 31'h253a_4255;
  assign p18_add_65274_comb = {p17_add_65170[1:0] ^ p17_add_65170[12:11] ^ p17_add_65170[21:20], p17_add_65170[31:21] ^ p17_add_65170[10:0] ^ p17_add_65170[19:9], p17_add_65170[20:12] ^ p17_add_65170[31:23] ^ p17_add_65170[8:0], p17_add_65170[11:2] ^ p17_add_65170[22:13] ^ p17_add_65170[31:22]} + (p18_and_65270_comb ^ p17_add_65170 & p17_add_64939 ^ p17_and_65165);
  assign p18_add_65251_comb = {p18_add_65224_comb[5:0] ^ p18_add_65224_comb[10:5] ^ p18_add_65224_comb[24:19], p18_add_65224_comb[31:27] ^ p18_add_65224_comb[4:0] ^ p18_add_65224_comb[18:14], p18_add_65224_comb[26:13] ^ p18_add_65224_comb[31:18] ^ p18_add_65224_comb[13:0], p18_add_65224_comb[12:6] ^ p18_add_65224_comb[17:11] ^ p18_add_65224_comb[31:25]} + p17_add_64892;
  assign p18_add_65252_comb = (p18_add_65224_comb & p17_add_65124 ^ ~(p18_add_65224_comb | ~p17_add_65020)) + {p18_add_65246_comb, p17_add_64411[0]};
  assign p18_add_65275_comb = p18_add_65223_comb + p18_add_65274_comb;
  assign p18_add_65253_comb = p18_add_65251_comb + p18_add_65252_comb;

  // Registers for pipe stage 18:
  reg [31:0] p18_add_65020;
  reg [31:0] p18_add_65124;
  reg [31:0] p18_add_65224;
  reg [31:0] p18_add_64939;
  reg [31:0] p18_add_65070;
  reg [31:0] p18_add_65170;
  reg [31:0] p18_and_65270;
  reg [31:0] p18_add_65275;
  reg [31:0] p18_add_64709;
  reg [31:0] p18_add_64264;
  reg [31:0] p18_add_64123;
  reg [31:0] p18_add_64692;
  reg [31:0] p18_add_64089;
  reg [31:0] p18_add_64569;
  reg [31:0] p18_add_64055;
  reg [31:0] p18_add_64551;
  reg [31:0] p18_add_64038;
  reg [31:0] p18_add_64429;
  reg [31:0] p18_add_64247;
  reg [31:0] p18_add_65253;
  reg [31:0] p18_add_64411;
  reg [31:0] p18_add_64001;
  reg [31:0] p18_add_63982;
  reg [31:0] p18_add_63945;
  reg [31:0] p18_add_63927;
  always_ff @ (posedge clk) begin
    p18_add_65020 <= p17_add_65020;
    p18_add_65124 <= p17_add_65124;
    p18_add_65224 <= p18_add_65224_comb;
    p18_add_64939 <= p17_add_64939;
    p18_add_65070 <= p17_add_65070;
    p18_add_65170 <= p17_add_65170;
    p18_and_65270 <= p18_and_65270_comb;
    p18_add_65275 <= p18_add_65275_comb;
    p18_add_64709 <= p17_add_64709;
    p18_add_64264 <= p17_add_64264;
    p18_add_64123 <= p17_add_64123;
    p18_add_64692 <= p17_add_64692;
    p18_add_64089 <= p17_add_64089;
    p18_add_64569 <= p17_add_64569;
    p18_add_64055 <= p17_add_64055;
    p18_add_64551 <= p17_add_64551;
    p18_add_64038 <= p17_add_64038;
    p18_add_64429 <= p17_add_64429;
    p18_add_64247 <= p17_add_64247;
    p18_add_65253 <= p18_add_65253_comb;
    p18_add_64411 <= p17_add_64411;
    p18_add_64001 <= p17_add_64001;
    p18_add_63982 <= p17_add_63982;
    p18_add_63945 <= p17_add_63945;
    p18_add_63927 <= p17_add_63927;
  end

  // ===== Pipe stage 19:
  wire [31:0] p19_and_65393_comb;
  wire [31:0] p19_add_65326_comb;
  wire [31:0] p19_add_65412_comb;
  wire [31:0] p19_add_65375_comb;
  wire [31:0] p19_add_65414_comb;
  wire [31:0] p19_add_65376_comb;
  wire [29:0] p19_add_65348_comb;
  wire [31:0] p19_and_65433_comb;
  wire [31:0] p19_add_65353_comb;
  wire [31:0] p19_add_65354_comb;
  wire [31:0] p19_add_65355_comb;
  wire [31:0] p19_add_65437_comb;
  wire [31:0] p19_add_65455_comb;
  wire [31:0] p19_add_65415_comb;
  wire [31:0] p19_add_65356_comb;
  wire [30:0] p19_add_65359_comb;
  wire [31:0] p19_add_65438_comb;
  wire [31:0] p19_add_65524_comb;
  wire [31:0] p19_add_65507_comb;
  wire [31:0] p19_add_65490_comb;
  wire [31:0] p19_add_65473_comb;
  wire [31:0] p19_add_65456_comb;
  wire [31:0] p19_add_65416_comb;
  assign p19_and_65393_comb = p18_add_65275 & p18_add_65170;
  assign p19_add_65326_comb = p18_add_64939 + p18_add_65253;
  assign p19_add_65412_comb = {p18_add_65275[1:0] ^ p18_add_65275[12:11] ^ p18_add_65275[21:20], p18_add_65275[31:21] ^ p18_add_65275[10:0] ^ p18_add_65275[19:9], p18_add_65275[20:12] ^ p18_add_65275[31:23] ^ p18_add_65275[8:0], p18_add_65275[11:2] ^ p18_add_65275[22:13] ^ p18_add_65275[31:22]} + (p19_and_65393_comb ^ p18_add_65275 & p18_add_65070 ^ p18_and_65270);
  assign p19_add_65375_comb = p18_add_63927 + {p18_add_64247[16:7] ^ p18_add_64247[18:9], p18_add_64247[6:0] ^ p18_add_64247[8:2] ^ p18_add_64247[31:25], p18_add_64247[31:30] ^ p18_add_64247[1:0] ^ p18_add_64247[24:23], p18_add_64247[29:17] ^ p18_add_64247[31:19] ^ p18_add_64247[22:10]};
  assign p19_add_65414_comb = p18_add_65253 + p19_add_65412_comb;
  assign p19_add_65376_comb = p18_add_64038 + p19_add_65375_comb;
  assign p19_add_65348_comb = p18_add_64247[31:2] + 30'h172c_2a77;
  assign p19_and_65433_comb = p19_add_65414_comb & p18_add_65275;
  assign p19_add_65353_comb = {p19_add_65326_comb[5:0] ^ p19_add_65326_comb[10:5] ^ p19_add_65326_comb[24:19], p19_add_65326_comb[31:27] ^ p19_add_65326_comb[4:0] ^ p19_add_65326_comb[18:14], p19_add_65326_comb[26:13] ^ p19_add_65326_comb[31:18] ^ p19_add_65326_comb[13:0], p19_add_65326_comb[12:6] ^ p19_add_65326_comb[17:11] ^ p19_add_65326_comb[31:25]} + p18_add_65020;
  assign p19_add_65354_comb = (p19_add_65326_comb & p18_add_65224 ^ ~(p19_add_65326_comb | ~p18_add_65124)) + {p19_add_65348_comb, p18_add_64247[1:0]};
  assign p19_add_65355_comb = p19_add_65353_comb + p19_add_65354_comb;
  assign p19_add_65437_comb = {p19_add_65414_comb[1:0] ^ p19_add_65414_comb[12:11] ^ p19_add_65414_comb[21:20], p19_add_65414_comb[31:21] ^ p19_add_65414_comb[10:0] ^ p19_add_65414_comb[19:9], p19_add_65414_comb[20:12] ^ p19_add_65414_comb[31:23] ^ p19_add_65414_comb[8:0], p19_add_65414_comb[11:2] ^ p19_add_65414_comb[22:13] ^ p19_add_65414_comb[31:22]} + (p19_and_65433_comb ^ p19_add_65414_comb & p18_add_65170 ^ p19_and_65393_comb);
  assign p19_add_65455_comb = p19_add_65376_comb + {p18_add_64692[16:7] ^ p18_add_64692[18:9], p18_add_64692[6:0] ^ p18_add_64692[8:2] ^ p18_add_64692[31:25], p18_add_64692[31:30] ^ p18_add_64692[1:0] ^ p18_add_64692[24:23], p18_add_64692[29:17] ^ p18_add_64692[31:19] ^ p18_add_64692[22:10]};
  assign p19_add_65415_comb = p18_add_63982 + {p19_add_65376_comb[16:7] ^ p19_add_65376_comb[18:9], p19_add_65376_comb[6:0] ^ p19_add_65376_comb[8:2] ^ p19_add_65376_comb[31:25], p19_add_65376_comb[31:30] ^ p19_add_65376_comb[1:0] ^ p19_add_65376_comb[24:23], p19_add_65376_comb[29:17] ^ p19_add_65376_comb[31:19] ^ p19_add_65376_comb[22:10]};
  assign p19_add_65356_comb = p18_add_65070 + p19_add_65355_comb;
  assign p19_add_65359_comb = p18_add_64429[31:1] + 31'h3b7c_c46d;
  assign p19_add_65438_comb = p19_add_65355_comb + p19_add_65437_comb;
  assign p19_add_65524_comb = {p18_add_64411[6:4] ^ p18_add_64411[17:15], p18_add_64411[3:0] ^ p18_add_64411[14:11] ^ p18_add_64411[31:28], p18_add_64411[31:21] ^ p18_add_64411[10:0] ^ p18_add_64411[27:17], p18_add_64411[20:7] ^ p18_add_64411[31:18] ^ p18_add_64411[16:3]} + p18_add_64001;
  assign p19_add_65507_comb = {p18_add_64001[6:4] ^ p18_add_64001[17:15], p18_add_64001[3:0] ^ p18_add_64001[14:11] ^ p18_add_64001[31:28], p18_add_64001[31:21] ^ p18_add_64001[10:0] ^ p18_add_64001[27:17], p18_add_64001[20:7] ^ p18_add_64001[31:18] ^ p18_add_64001[16:3]} + p18_add_63982;
  assign p19_add_65490_comb = {p18_add_63982[6:4] ^ p18_add_63982[17:15], p18_add_63982[3:0] ^ p18_add_63982[14:11] ^ p18_add_63982[31:28], p18_add_63982[31:21] ^ p18_add_63982[10:0] ^ p18_add_63982[27:17], p18_add_63982[20:7] ^ p18_add_63982[31:18] ^ p18_add_63982[16:3]} + p18_add_63945;
  assign p19_add_65473_comb = {p18_add_63945[6:4] ^ p18_add_63945[17:15], p18_add_63945[3:0] ^ p18_add_63945[14:11] ^ p18_add_63945[31:28], p18_add_63945[31:21] ^ p18_add_63945[10:0] ^ p18_add_63945[27:17], p18_add_63945[20:7] ^ p18_add_63945[31:18] ^ p18_add_63945[16:3]} + p18_add_63927;
  assign p19_add_65456_comb = p18_add_64264 + p19_add_65455_comb;
  assign p19_add_65416_comb = p18_add_64055 + p19_add_65415_comb;

  // Registers for pipe stage 19:
  reg [31:0] p19_add_65124;
  reg [31:0] p19_add_65224;
  reg [31:0] p19_add_65326;
  reg [31:0] p19_add_65356;
  reg [30:0] p19_add_65359;
  reg [31:0] p19_add_65170;
  reg [31:0] p19_add_65275;
  reg [31:0] p19_add_65414;
  reg [31:0] p19_and_65433;
  reg [31:0] p19_add_65438;
  reg [31:0] p19_add_65524;
  reg [31:0] p19_add_65507;
  reg [31:0] p19_add_65490;
  reg [31:0] p19_add_65473;
  reg [31:0] p19_add_64709;
  reg [31:0] p19_add_65456;
  reg [31:0] p19_add_64123;
  reg [31:0] p19_add_64692;
  reg [31:0] p19_add_64089;
  reg [31:0] p19_add_64569;
  reg [31:0] p19_add_65416;
  reg [31:0] p19_add_64551;
  reg [31:0] p19_add_65376;
  reg [31:0] p19_add_64429;
  reg [31:0] p19_add_64247;
  reg [31:0] p19_add_64411;
  always_ff @ (posedge clk) begin
    p19_add_65124 <= p18_add_65124;
    p19_add_65224 <= p18_add_65224;
    p19_add_65326 <= p19_add_65326_comb;
    p19_add_65356 <= p19_add_65356_comb;
    p19_add_65359 <= p19_add_65359_comb;
    p19_add_65170 <= p18_add_65170;
    p19_add_65275 <= p18_add_65275;
    p19_add_65414 <= p19_add_65414_comb;
    p19_and_65433 <= p19_and_65433_comb;
    p19_add_65438 <= p19_add_65438_comb;
    p19_add_65524 <= p19_add_65524_comb;
    p19_add_65507 <= p19_add_65507_comb;
    p19_add_65490 <= p19_add_65490_comb;
    p19_add_65473 <= p19_add_65473_comb;
    p19_add_64709 <= p18_add_64709;
    p19_add_65456 <= p19_add_65456_comb;
    p19_add_64123 <= p18_add_64123;
    p19_add_64692 <= p18_add_64692;
    p19_add_64089 <= p18_add_64089;
    p19_add_64569 <= p18_add_64569;
    p19_add_65416 <= p19_add_65416_comb;
    p19_add_64551 <= p18_add_64551;
    p19_add_65376 <= p19_add_65376_comb;
    p19_add_64429 <= p18_add_64429;
    p19_add_64247 <= p18_add_64247;
    p19_add_64411 <= p18_add_64411;
  end

  // ===== Pipe stage 20:
  wire [31:0] p20_add_65707_comb;
  wire [31:0] p20_add_65671_comb;
  wire [31:0] p20_add_65600_comb;
  wire [31:0] p20_add_65601_comb;
  wire [31:0] p20_add_65708_comb;
  wire [31:0] p20_add_65672_comb;
  wire [31:0] p20_add_65602_comb;
  wire [31:0] p20_add_65603_comb;
  wire [31:0] p20_and_65649_comb;
  wire [30:0] p20_add_65625_comb;
  wire [31:0] p20_add_65653_comb;
  wire [31:0] p20_add_65725_comb;
  wire [31:0] p20_add_65689_comb;
  wire [31:0] p20_add_65632_comb;
  wire [31:0] p20_add_65654_comb;
  wire [31:0] p20_add_65794_comb;
  wire [31:0] p20_add_65777_comb;
  wire [31:0] p20_add_65760_comb;
  wire [31:0] p20_add_65743_comb;
  wire [31:0] p20_add_65726_comb;
  wire [31:0] p20_add_65690_comb;
  wire [31:0] p20_add_65630_comb;
  wire [31:0] p20_add_65631_comb;
  assign p20_add_65707_comb = p19_add_65416 + {p19_add_65456[16:7] ^ p19_add_65456[18:9], p19_add_65456[6:0] ^ p19_add_65456[8:2] ^ p19_add_65456[31:25], p19_add_65456[31:30] ^ p19_add_65456[1:0] ^ p19_add_65456[24:23], p19_add_65456[29:17] ^ p19_add_65456[31:19] ^ p19_add_65456[22:10]};
  assign p20_add_65671_comb = p19_add_64411 + {p19_add_65416[16:7] ^ p19_add_65416[18:9], p19_add_65416[6:0] ^ p19_add_65416[8:2] ^ p19_add_65416[31:25], p19_add_65416[31:30] ^ p19_add_65416[1:0] ^ p19_add_65416[24:23], p19_add_65416[29:17] ^ p19_add_65416[31:19] ^ p19_add_65416[22:10]};
  assign p20_add_65600_comb = {p19_add_65356[5:0] ^ p19_add_65356[10:5] ^ p19_add_65356[24:19], p19_add_65356[31:27] ^ p19_add_65356[4:0] ^ p19_add_65356[18:14], p19_add_65356[26:13] ^ p19_add_65356[31:18] ^ p19_add_65356[13:0], p19_add_65356[12:6] ^ p19_add_65356[17:11] ^ p19_add_65356[31:25]} + p19_add_65124;
  assign p20_add_65601_comb = (p19_add_65356 & p19_add_65326 ^ ~(p19_add_65356 | ~p19_add_65224)) + {p19_add_65359, p19_add_64429[0]};
  assign p20_add_65708_comb = p19_add_65473 + p20_add_65707_comb;
  assign p20_add_65672_comb = p19_add_64089 + p20_add_65671_comb;
  assign p20_add_65602_comb = p20_add_65600_comb + p20_add_65601_comb;
  assign p20_add_65603_comb = p19_add_65170 + p20_add_65602_comb;
  assign p20_and_65649_comb = p19_add_65438 & p19_add_65414;
  assign p20_add_65625_comb = p19_add_65376[31:1] + 31'h4c1f_28a9;
  assign p20_add_65653_comb = {p19_add_65438[1:0] ^ p19_add_65438[12:11] ^ p19_add_65438[21:20], p19_add_65438[31:21] ^ p19_add_65438[10:0] ^ p19_add_65438[19:9], p19_add_65438[20:12] ^ p19_add_65438[31:23] ^ p19_add_65438[8:0], p19_add_65438[11:2] ^ p19_add_65438[22:13] ^ p19_add_65438[31:22]} + (p20_and_65649_comb ^ p19_add_65438 & p19_add_65275 ^ p19_and_65433);
  assign p20_add_65725_comb = p20_add_65672_comb + {p20_add_65708_comb[16:7] ^ p20_add_65708_comb[18:9], p20_add_65708_comb[6:0] ^ p20_add_65708_comb[8:2] ^ p20_add_65708_comb[31:25], p20_add_65708_comb[31:30] ^ p20_add_65708_comb[1:0] ^ p20_add_65708_comb[24:23], p20_add_65708_comb[29:17] ^ p20_add_65708_comb[31:19] ^ p20_add_65708_comb[22:10]};
  assign p20_add_65689_comb = p19_add_64429 + {p20_add_65672_comb[16:7] ^ p20_add_65672_comb[18:9], p20_add_65672_comb[6:0] ^ p20_add_65672_comb[8:2] ^ p20_add_65672_comb[31:25], p20_add_65672_comb[31:30] ^ p20_add_65672_comb[1:0] ^ p20_add_65672_comb[24:23], p20_add_65672_comb[29:17] ^ p20_add_65672_comb[31:19] ^ p20_add_65672_comb[22:10]};
  assign p20_add_65632_comb = p19_add_65326 + p19_add_64551;
  assign p20_add_65654_comb = p20_add_65602_comb + p20_add_65653_comb;
  assign p20_add_65794_comb = {p19_add_64551[6:4] ^ p19_add_64551[17:15], p19_add_64551[3:0] ^ p19_add_64551[14:11] ^ p19_add_64551[31:28], p19_add_64551[31:21] ^ p19_add_64551[10:0] ^ p19_add_64551[27:17], p19_add_64551[20:7] ^ p19_add_64551[31:18] ^ p19_add_64551[16:3]} + p19_add_65376;
  assign p20_add_65777_comb = {p19_add_65376[6:4] ^ p19_add_65376[17:15], p19_add_65376[3:0] ^ p19_add_65376[14:11] ^ p19_add_65376[31:28], p19_add_65376[31:21] ^ p19_add_65376[10:0] ^ p19_add_65376[27:17], p19_add_65376[20:7] ^ p19_add_65376[31:18] ^ p19_add_65376[16:3]} + p19_add_64429;
  assign p20_add_65760_comb = {p19_add_64429[6:4] ^ p19_add_64429[17:15], p19_add_64429[3:0] ^ p19_add_64429[14:11] ^ p19_add_64429[31:28], p19_add_64429[31:21] ^ p19_add_64429[10:0] ^ p19_add_64429[27:17], p19_add_64429[20:7] ^ p19_add_64429[31:18] ^ p19_add_64429[16:3]} + p19_add_64247;
  assign p20_add_65743_comb = {p19_add_64247[6:4] ^ p19_add_64247[17:15], p19_add_64247[3:0] ^ p19_add_64247[14:11] ^ p19_add_64247[31:28], p19_add_64247[31:21] ^ p19_add_64247[10:0] ^ p19_add_64247[27:17], p19_add_64247[20:7] ^ p19_add_64247[31:18] ^ p19_add_64247[16:3]} + p19_add_64411;
  assign p20_add_65726_comb = p19_add_65507 + p20_add_65725_comb;
  assign p20_add_65690_comb = p19_add_64123 + p20_add_65689_comb;
  assign p20_add_65630_comb = {p20_add_65603_comb[5:0] ^ p20_add_65603_comb[10:5] ^ p20_add_65603_comb[24:19], p20_add_65603_comb[31:27] ^ p20_add_65603_comb[4:0] ^ p20_add_65603_comb[18:14], p20_add_65603_comb[26:13] ^ p20_add_65603_comb[31:18] ^ p20_add_65603_comb[13:0], p20_add_65603_comb[12:6] ^ p20_add_65603_comb[17:11] ^ p20_add_65603_comb[31:25]} + p19_add_65224;
  assign p20_add_65631_comb = (p20_add_65603_comb & p19_add_65356 ^ ~(p20_add_65603_comb | ~p19_add_65326)) + {p20_add_65625_comb, p19_add_65376[0]};

  // Registers for pipe stage 20:
  reg [31:0] p20_add_65356;
  reg [31:0] p20_add_65603;
  reg [31:0] p20_add_65275;
  reg [31:0] p20_add_65632;
  reg [31:0] p20_add_65414;
  reg [31:0] p20_add_65438;
  reg [31:0] p20_and_65649;
  reg [31:0] p20_add_65654;
  reg [31:0] p20_add_65794;
  reg [31:0] p20_add_65777;
  reg [31:0] p20_add_65760;
  reg [31:0] p20_add_65743;
  reg [31:0] p20_add_65524;
  reg [31:0] p20_add_65726;
  reg [31:0] p20_add_65490;
  reg [31:0] p20_add_65708;
  reg [31:0] p20_add_64709;
  reg [31:0] p20_add_65456;
  reg [31:0] p20_add_65690;
  reg [31:0] p20_add_64692;
  reg [31:0] p20_add_65672;
  reg [31:0] p20_add_64569;
  reg [31:0] p20_add_65416;
  reg [31:0] p20_add_64551;
  reg [31:0] p20_add_65630;
  reg [31:0] p20_add_65631;
  always_ff @ (posedge clk) begin
    p20_add_65356 <= p19_add_65356;
    p20_add_65603 <= p20_add_65603_comb;
    p20_add_65275 <= p19_add_65275;
    p20_add_65632 <= p20_add_65632_comb;
    p20_add_65414 <= p19_add_65414;
    p20_add_65438 <= p19_add_65438;
    p20_and_65649 <= p20_and_65649_comb;
    p20_add_65654 <= p20_add_65654_comb;
    p20_add_65794 <= p20_add_65794_comb;
    p20_add_65777 <= p20_add_65777_comb;
    p20_add_65760 <= p20_add_65760_comb;
    p20_add_65743 <= p20_add_65743_comb;
    p20_add_65524 <= p19_add_65524;
    p20_add_65726 <= p20_add_65726_comb;
    p20_add_65490 <= p19_add_65490;
    p20_add_65708 <= p20_add_65708_comb;
    p20_add_64709 <= p19_add_64709;
    p20_add_65456 <= p19_add_65456;
    p20_add_65690 <= p20_add_65690_comb;
    p20_add_64692 <= p19_add_64692;
    p20_add_65672 <= p20_add_65672_comb;
    p20_add_64569 <= p19_add_64569;
    p20_add_65416 <= p19_add_65416;
    p20_add_64551 <= p19_add_64551;
    p20_add_65630 <= p20_add_65630_comb;
    p20_add_65631 <= p20_add_65631_comb;
  end

  // ===== Pipe stage 21:
  wire [31:0] p21_add_65847_comb;
  wire [31:0] p21_add_65947_comb;
  wire [31:0] p21_add_65911_comb;
  wire [31:0] p21_add_65848_comb;
  wire [31:0] p21_add_65948_comb;
  wire [31:0] p21_add_65912_comb;
  wire [31:0] p21_and_65889_comb;
  wire [31:0] p21_add_65893_comb;
  wire [31:0] p21_add_65870_comb;
  wire [31:0] p21_add_65965_comb;
  wire [31:0] p21_add_65929_comb;
  wire [31:0] p21_add_65894_comb;
  wire [31:0] p21_add_65872_comb;
  wire [31:0] p21_add_65983_comb;
  wire [31:0] p21_add_65966_comb;
  wire [31:0] p21_add_65930_comb;
  assign p21_add_65847_comb = p20_add_65630 + p20_add_65631;
  assign p21_add_65947_comb = p20_add_65690 + {p20_add_65726[16:7] ^ p20_add_65726[18:9], p20_add_65726[6:0] ^ p20_add_65726[8:2] ^ p20_add_65726[31:25], p20_add_65726[31:30] ^ p20_add_65726[1:0] ^ p20_add_65726[24:23], p20_add_65726[29:17] ^ p20_add_65726[31:19] ^ p20_add_65726[22:10]};
  assign p21_add_65911_comb = p20_add_64551 + {p20_add_65690[16:7] ^ p20_add_65690[18:9], p20_add_65690[6:0] ^ p20_add_65690[8:2] ^ p20_add_65690[31:25], p20_add_65690[31:30] ^ p20_add_65690[1:0] ^ p20_add_65690[24:23], p20_add_65690[29:17] ^ p20_add_65690[31:19] ^ p20_add_65690[22:10]};
  assign p21_add_65848_comb = p20_add_65275 + p21_add_65847_comb;
  assign p21_add_65948_comb = p20_add_65743 + p21_add_65947_comb;
  assign p21_add_65912_comb = p20_add_64709 + p21_add_65911_comb;
  assign p21_and_65889_comb = p20_add_65654 & p20_add_65438;
  assign p21_add_65893_comb = {p20_add_65654[1:0] ^ p20_add_65654[12:11] ^ p20_add_65654[21:20], p20_add_65654[31:21] ^ p20_add_65654[10:0] ^ p20_add_65654[19:9], p20_add_65654[20:12] ^ p20_add_65654[31:23] ^ p20_add_65654[8:0], p20_add_65654[11:2] ^ p20_add_65654[22:13] ^ p20_add_65654[31:22]} + (p21_and_65889_comb ^ p20_add_65654 & p20_add_65414 ^ p20_and_65649);
  assign p21_add_65870_comb = {p21_add_65848_comb[5:0] ^ p21_add_65848_comb[10:5] ^ p21_add_65848_comb[24:19], p21_add_65848_comb[31:27] ^ p21_add_65848_comb[4:0] ^ p21_add_65848_comb[18:14], p21_add_65848_comb[26:13] ^ p21_add_65848_comb[31:18] ^ p21_add_65848_comb[13:0], p21_add_65848_comb[12:6] ^ p21_add_65848_comb[17:11] ^ p21_add_65848_comb[31:25]} + (p21_add_65848_comb & p20_add_65603 ^ ~(p21_add_65848_comb | ~p20_add_65356));
  assign p21_add_65965_comb = p21_add_65912_comb + {p21_add_65948_comb[16:7] ^ p21_add_65948_comb[18:9], p21_add_65948_comb[6:0] ^ p21_add_65948_comb[8:2] ^ p21_add_65948_comb[31:25], p21_add_65948_comb[31:30] ^ p21_add_65948_comb[1:0] ^ p21_add_65948_comb[24:23], p21_add_65948_comb[29:17] ^ p21_add_65948_comb[31:19] ^ p21_add_65948_comb[22:10]};
  assign p21_add_65929_comb = p20_add_64569 + {p21_add_65912_comb[16:7] ^ p21_add_65912_comb[18:9], p21_add_65912_comb[6:0] ^ p21_add_65912_comb[8:2] ^ p21_add_65912_comb[31:25], p21_add_65912_comb[31:30] ^ p21_add_65912_comb[1:0] ^ p21_add_65912_comb[24:23], p21_add_65912_comb[29:17] ^ p21_add_65912_comb[31:19] ^ p21_add_65912_comb[22:10]};
  assign p21_add_65894_comb = p21_add_65847_comb + p21_add_65893_comb;
  assign p21_add_65872_comb = p21_add_65870_comb + 32'ha831_c66d;
  assign p21_add_65983_comb = {p20_add_65416[6:4] ^ p20_add_65416[17:15], p20_add_65416[3:0] ^ p20_add_65416[14:11] ^ p20_add_65416[31:28], p20_add_65416[31:21] ^ p20_add_65416[10:0] ^ p20_add_65416[27:17], p20_add_65416[20:7] ^ p20_add_65416[31:18] ^ p20_add_65416[16:3]} + p20_add_64551;
  assign p21_add_65966_comb = p20_add_65777 + p21_add_65965_comb;
  assign p21_add_65930_comb = p20_add_65490 + p21_add_65929_comb;

  // Registers for pipe stage 21:
  reg [31:0] p21_add_65356;
  reg [31:0] p21_add_65603;
  reg [31:0] p21_add_65848;
  reg [31:0] p21_add_65632;
  reg [31:0] p21_add_65414;
  reg [31:0] p21_add_65438;
  reg [31:0] p21_add_65654;
  reg [31:0] p21_and_65889;
  reg [31:0] p21_add_65894;
  reg [31:0] p21_add_65872;
  reg [31:0] p21_add_65983;
  reg [31:0] p21_add_65794;
  reg [31:0] p21_add_65966;
  reg [31:0] p21_add_65760;
  reg [31:0] p21_add_65948;
  reg [31:0] p21_add_65524;
  reg [31:0] p21_add_65726;
  reg [31:0] p21_add_65930;
  reg [31:0] p21_add_65708;
  reg [31:0] p21_add_65912;
  reg [31:0] p21_add_65456;
  reg [31:0] p21_add_65690;
  reg [31:0] p21_add_64692;
  reg [31:0] p21_add_65672;
  reg [31:0] p21_add_64569;
  reg [31:0] p21_add_65416;
  always_ff @ (posedge clk) begin
    p21_add_65356 <= p20_add_65356;
    p21_add_65603 <= p20_add_65603;
    p21_add_65848 <= p21_add_65848_comb;
    p21_add_65632 <= p20_add_65632;
    p21_add_65414 <= p20_add_65414;
    p21_add_65438 <= p20_add_65438;
    p21_add_65654 <= p20_add_65654;
    p21_and_65889 <= p21_and_65889_comb;
    p21_add_65894 <= p21_add_65894_comb;
    p21_add_65872 <= p21_add_65872_comb;
    p21_add_65983 <= p21_add_65983_comb;
    p21_add_65794 <= p20_add_65794;
    p21_add_65966 <= p21_add_65966_comb;
    p21_add_65760 <= p20_add_65760;
    p21_add_65948 <= p21_add_65948_comb;
    p21_add_65524 <= p20_add_65524;
    p21_add_65726 <= p20_add_65726;
    p21_add_65930 <= p21_add_65930_comb;
    p21_add_65708 <= p20_add_65708;
    p21_add_65912 <= p21_add_65912_comb;
    p21_add_65456 <= p20_add_65456;
    p21_add_65690 <= p20_add_65690;
    p21_add_64692 <= p20_add_64692;
    p21_add_65672 <= p20_add_65672;
    p21_add_64569 <= p20_add_64569;
    p21_add_65416 <= p20_add_65416;
  end

  // ===== Pipe stage 22:
  wire [31:0] p22_add_66036_comb;
  wire [31:0] p22_add_66037_comb;
  wire [31:0] p22_and_66084_comb;
  wire [28:0] p22_add_66059_comb;
  wire [31:0] p22_add_66088_comb;
  wire [31:0] p22_add_66106_comb;
  wire [31:0] p22_add_66064_comb;
  wire [31:0] p22_add_66065_comb;
  wire [31:0] p22_add_66067_comb;
  wire [31:0] p22_add_66089_comb;
  wire [31:0] p22_add_66141_comb;
  wire [31:0] p22_add_66124_comb;
  wire [31:0] p22_add_66118_comb;
  wire [31:0] p22_add_66066_comb;
  assign p22_add_66036_comb = p21_add_65872 + p21_add_65632;
  assign p22_add_66037_comb = p21_add_65414 + p22_add_66036_comb;
  assign p22_and_66084_comb = p21_add_65894 & p21_add_65654;
  assign p22_add_66059_comb = p21_add_65416[31:3] + 29'h1600_64f9;
  assign p22_add_66088_comb = {p21_add_65894[1:0] ^ p21_add_65894[12:11] ^ p21_add_65894[21:20], p21_add_65894[31:21] ^ p21_add_65894[10:0] ^ p21_add_65894[19:9], p21_add_65894[20:12] ^ p21_add_65894[31:23] ^ p21_add_65894[8:0], p21_add_65894[11:2] ^ p21_add_65894[22:13] ^ p21_add_65894[31:22]} + (p22_and_66084_comb ^ p21_add_65894 & p21_add_65438 ^ p21_and_65889);
  assign p22_add_66106_comb = p21_add_65930 + {p21_add_65966[16:7] ^ p21_add_65966[18:9], p21_add_65966[6:0] ^ p21_add_65966[8:2] ^ p21_add_65966[31:25], p21_add_65966[31:30] ^ p21_add_65966[1:0] ^ p21_add_65966[24:23], p21_add_65966[29:17] ^ p21_add_65966[31:19] ^ p21_add_65966[22:10]};
  assign p22_add_66064_comb = {p22_add_66037_comb[5:0] ^ p22_add_66037_comb[10:5] ^ p22_add_66037_comb[24:19], p22_add_66037_comb[31:27] ^ p22_add_66037_comb[4:0] ^ p22_add_66037_comb[18:14], p22_add_66037_comb[26:13] ^ p22_add_66037_comb[31:18] ^ p22_add_66037_comb[13:0], p22_add_66037_comb[12:6] ^ p22_add_66037_comb[17:11] ^ p22_add_66037_comb[31:25]} + p21_add_65356;
  assign p22_add_66065_comb = (p22_add_66037_comb & p21_add_65848 ^ ~(p22_add_66037_comb | ~p21_add_65603)) + {p22_add_66059_comb, p21_add_65416[2:0]};
  assign p22_add_66067_comb = p21_add_65603 + p21_add_64569;
  assign p22_add_66089_comb = p22_add_66036_comb + p22_add_66088_comb;
  assign p22_add_66141_comb = {p21_add_65672[6:4] ^ p21_add_65672[17:15], p21_add_65672[3:0] ^ p21_add_65672[14:11] ^ p21_add_65672[31:28], p21_add_65672[31:21] ^ p21_add_65672[10:0] ^ p21_add_65672[27:17], p21_add_65672[20:7] ^ p21_add_65672[31:18] ^ p21_add_65672[16:3]} + p21_add_64569;
  assign p22_add_66124_comb = {p21_add_64569[6:4] ^ p21_add_64569[17:15], p21_add_64569[3:0] ^ p21_add_64569[14:11] ^ p21_add_64569[31:28], p21_add_64569[31:21] ^ p21_add_64569[10:0] ^ p21_add_64569[27:17], p21_add_64569[20:7] ^ p21_add_64569[31:18] ^ p21_add_64569[16:3]} + p21_add_65416;
  assign p22_add_66118_comb = p21_add_65983 + p22_add_66106_comb;
  assign p22_add_66066_comb = p22_add_66064_comb + p22_add_66065_comb;

  // Registers for pipe stage 22:
  reg [31:0] p22_add_65848;
  reg [31:0] p22_add_66037;
  reg [31:0] p22_add_65438;
  reg [31:0] p22_add_66067;
  reg [31:0] p22_add_65654;
  reg [31:0] p22_add_65894;
  reg [31:0] p22_and_66084;
  reg [31:0] p22_add_66089;
  reg [31:0] p22_add_66141;
  reg [31:0] p22_add_66124;
  reg [31:0] p22_add_66118;
  reg [31:0] p22_add_65794;
  reg [31:0] p22_add_65966;
  reg [31:0] p22_add_65760;
  reg [31:0] p22_add_65948;
  reg [31:0] p22_add_65524;
  reg [31:0] p22_add_65726;
  reg [31:0] p22_add_65930;
  reg [31:0] p22_add_65708;
  reg [31:0] p22_add_65912;
  reg [31:0] p22_add_65456;
  reg [31:0] p22_add_65690;
  reg [31:0] p22_add_64692;
  reg [31:0] p22_add_65672;
  reg [31:0] p22_add_66066;
  always_ff @ (posedge clk) begin
    p22_add_65848 <= p21_add_65848;
    p22_add_66037 <= p22_add_66037_comb;
    p22_add_65438 <= p21_add_65438;
    p22_add_66067 <= p22_add_66067_comb;
    p22_add_65654 <= p21_add_65654;
    p22_add_65894 <= p21_add_65894;
    p22_and_66084 <= p22_and_66084_comb;
    p22_add_66089 <= p22_add_66089_comb;
    p22_add_66141 <= p22_add_66141_comb;
    p22_add_66124 <= p22_add_66124_comb;
    p22_add_66118 <= p22_add_66118_comb;
    p22_add_65794 <= p21_add_65794;
    p22_add_65966 <= p21_add_65966;
    p22_add_65760 <= p21_add_65760;
    p22_add_65948 <= p21_add_65948;
    p22_add_65524 <= p21_add_65524;
    p22_add_65726 <= p21_add_65726;
    p22_add_65930 <= p21_add_65930;
    p22_add_65708 <= p21_add_65708;
    p22_add_65912 <= p21_add_65912;
    p22_add_65456 <= p21_add_65456;
    p22_add_65690 <= p21_add_65690;
    p22_add_64692 <= p21_add_64692;
    p22_add_65672 <= p21_add_65672;
    p22_add_66066 <= p22_add_66066_comb;
  end

  // ===== Pipe stage 23:
  wire [31:0] p23_add_66192_comb;
  wire [31:0] p23_and_66235_comb;
  wire [31:0] p23_add_66214_comb;
  wire [31:0] p23_add_66216_comb;
  wire [31:0] p23_add_66239_comb;
  wire [31:0] p23_add_66217_comb;
  wire [31:0] p23_add_66218_comb;
  wire [31:0] p23_add_66240_comb;
  wire [31:0] p23_add_66257_comb;
  assign p23_add_66192_comb = p22_add_65438 + p22_add_66066;
  assign p23_and_66235_comb = p22_add_66089 & p22_add_65894;
  assign p23_add_66214_comb = {p23_add_66192_comb[5:0] ^ p23_add_66192_comb[10:5] ^ p23_add_66192_comb[24:19], p23_add_66192_comb[31:27] ^ p23_add_66192_comb[4:0] ^ p23_add_66192_comb[18:14], p23_add_66192_comb[26:13] ^ p23_add_66192_comb[31:18] ^ p23_add_66192_comb[13:0], p23_add_66192_comb[12:6] ^ p23_add_66192_comb[17:11] ^ p23_add_66192_comb[31:25]} + (p23_add_66192_comb & p22_add_66037 ^ ~(p23_add_66192_comb | ~p22_add_65848));
  assign p23_add_66216_comb = p23_add_66214_comb + 32'hbf59_7fc7;
  assign p23_add_66239_comb = {p22_add_66089[1:0] ^ p22_add_66089[12:11] ^ p22_add_66089[21:20], p22_add_66089[31:21] ^ p22_add_66089[10:0] ^ p22_add_66089[19:9], p22_add_66089[20:12] ^ p22_add_66089[31:23] ^ p22_add_66089[8:0], p22_add_66089[11:2] ^ p22_add_66089[22:13] ^ p22_add_66089[31:22]} + (p23_and_66235_comb ^ p22_add_66089 & p22_add_65654 ^ p22_and_66084);
  assign p23_add_66217_comb = p23_add_66216_comb + p22_add_66067;
  assign p23_add_66218_comb = p22_add_65848 + p22_add_65672;
  assign p23_add_66240_comb = p22_add_66066 + p23_add_66239_comb;
  assign p23_add_66257_comb = {p22_add_64692[6:4] ^ p22_add_64692[17:15], p22_add_64692[3:0] ^ p22_add_64692[14:11] ^ p22_add_64692[31:28], p22_add_64692[31:21] ^ p22_add_64692[10:0] ^ p22_add_64692[27:17], p22_add_64692[20:7] ^ p22_add_64692[31:18] ^ p22_add_64692[16:3]} + p22_add_65672;

  // Registers for pipe stage 23:
  reg [31:0] p23_add_66037;
  reg [31:0] p23_add_66192;
  reg [31:0] p23_add_65654;
  reg [31:0] p23_add_66217;
  reg [31:0] p23_add_66218;
  reg [31:0] p23_add_65894;
  reg [31:0] p23_add_66089;
  reg [31:0] p23_and_66235;
  reg [31:0] p23_add_66240;
  reg [31:0] p23_add_66257;
  reg [31:0] p23_add_66141;
  reg [31:0] p23_add_66124;
  reg [31:0] p23_add_66118;
  reg [31:0] p23_add_65794;
  reg [31:0] p23_add_65966;
  reg [31:0] p23_add_65760;
  reg [31:0] p23_add_65948;
  reg [31:0] p23_add_65524;
  reg [31:0] p23_add_65726;
  reg [31:0] p23_add_65930;
  reg [31:0] p23_add_65708;
  reg [31:0] p23_add_65912;
  reg [31:0] p23_add_65456;
  reg [31:0] p23_add_65690;
  reg [31:0] p23_add_64692;
  always_ff @ (posedge clk) begin
    p23_add_66037 <= p22_add_66037;
    p23_add_66192 <= p23_add_66192_comb;
    p23_add_65654 <= p22_add_65654;
    p23_add_66217 <= p23_add_66217_comb;
    p23_add_66218 <= p23_add_66218_comb;
    p23_add_65894 <= p22_add_65894;
    p23_add_66089 <= p22_add_66089;
    p23_and_66235 <= p23_and_66235_comb;
    p23_add_66240 <= p23_add_66240_comb;
    p23_add_66257 <= p23_add_66257_comb;
    p23_add_66141 <= p22_add_66141;
    p23_add_66124 <= p22_add_66124;
    p23_add_66118 <= p22_add_66118;
    p23_add_65794 <= p22_add_65794;
    p23_add_65966 <= p22_add_65966;
    p23_add_65760 <= p22_add_65760;
    p23_add_65948 <= p22_add_65948;
    p23_add_65524 <= p22_add_65524;
    p23_add_65726 <= p22_add_65726;
    p23_add_65930 <= p22_add_65930;
    p23_add_65708 <= p22_add_65708;
    p23_add_65912 <= p22_add_65912;
    p23_add_65456 <= p22_add_65456;
    p23_add_65690 <= p22_add_65690;
    p23_add_64692 <= p22_add_64692;
  end

  // ===== Pipe stage 24:
  wire [31:0] p24_add_66308_comb;
  wire [31:0] p24_and_66351_comb;
  wire [31:0] p24_add_66330_comb;
  wire [31:0] p24_add_66332_comb;
  wire [31:0] p24_add_66355_comb;
  wire [31:0] p24_add_66333_comb;
  wire [31:0] p24_add_66334_comb;
  wire [31:0] p24_add_66356_comb;
  assign p24_add_66308_comb = p23_add_65654 + p23_add_66217;
  assign p24_and_66351_comb = p23_add_66240 & p23_add_66089;
  assign p24_add_66330_comb = {p24_add_66308_comb[5:0] ^ p24_add_66308_comb[10:5] ^ p24_add_66308_comb[24:19], p24_add_66308_comb[31:27] ^ p24_add_66308_comb[4:0] ^ p24_add_66308_comb[18:14], p24_add_66308_comb[26:13] ^ p24_add_66308_comb[31:18] ^ p24_add_66308_comb[13:0], p24_add_66308_comb[12:6] ^ p24_add_66308_comb[17:11] ^ p24_add_66308_comb[31:25]} + (p24_add_66308_comb & p23_add_66192 ^ ~(p24_add_66308_comb | ~p23_add_66037));
  assign p24_add_66332_comb = p24_add_66330_comb + 32'hc6e0_0bf3;
  assign p24_add_66355_comb = {p23_add_66240[1:0] ^ p23_add_66240[12:11] ^ p23_add_66240[21:20], p23_add_66240[31:21] ^ p23_add_66240[10:0] ^ p23_add_66240[19:9], p23_add_66240[20:12] ^ p23_add_66240[31:23] ^ p23_add_66240[8:0], p23_add_66240[11:2] ^ p23_add_66240[22:13] ^ p23_add_66240[31:22]} + (p24_and_66351_comb ^ p23_add_66240 & p23_add_65894 ^ p23_and_66235);
  assign p24_add_66333_comb = p24_add_66332_comb + p23_add_66218;
  assign p24_add_66334_comb = p23_add_66037 + p23_add_64692;
  assign p24_add_66356_comb = p23_add_66217 + p24_add_66355_comb;

  // Registers for pipe stage 24:
  reg [31:0] p24_add_66192;
  reg [31:0] p24_add_66308;
  reg [31:0] p24_add_65894;
  reg [31:0] p24_add_66333;
  reg [31:0] p24_add_66334;
  reg [31:0] p24_add_66089;
  reg [31:0] p24_add_66240;
  reg [31:0] p24_and_66351;
  reg [31:0] p24_add_66356;
  reg [31:0] p24_add_66257;
  reg [31:0] p24_add_66141;
  reg [31:0] p24_add_66124;
  reg [31:0] p24_add_66118;
  reg [31:0] p24_add_65794;
  reg [31:0] p24_add_65966;
  reg [31:0] p24_add_65760;
  reg [31:0] p24_add_65948;
  reg [31:0] p24_add_65524;
  reg [31:0] p24_add_65726;
  reg [31:0] p24_add_65930;
  reg [31:0] p24_add_65708;
  reg [31:0] p24_add_65912;
  reg [31:0] p24_add_65456;
  reg [31:0] p24_add_65690;
  reg [31:0] p24_add_64692;
  always_ff @ (posedge clk) begin
    p24_add_66192 <= p23_add_66192;
    p24_add_66308 <= p24_add_66308_comb;
    p24_add_65894 <= p23_add_65894;
    p24_add_66333 <= p24_add_66333_comb;
    p24_add_66334 <= p24_add_66334_comb;
    p24_add_66089 <= p23_add_66089;
    p24_add_66240 <= p23_add_66240;
    p24_and_66351 <= p24_and_66351_comb;
    p24_add_66356 <= p24_add_66356_comb;
    p24_add_66257 <= p23_add_66257;
    p24_add_66141 <= p23_add_66141;
    p24_add_66124 <= p23_add_66124;
    p24_add_66118 <= p23_add_66118;
    p24_add_65794 <= p23_add_65794;
    p24_add_65966 <= p23_add_65966;
    p24_add_65760 <= p23_add_65760;
    p24_add_65948 <= p23_add_65948;
    p24_add_65524 <= p23_add_65524;
    p24_add_65726 <= p23_add_65726;
    p24_add_65930 <= p23_add_65930;
    p24_add_65708 <= p23_add_65708;
    p24_add_65912 <= p23_add_65912;
    p24_add_65456 <= p23_add_65456;
    p24_add_65690 <= p23_add_65690;
    p24_add_64692 <= p23_add_64692;
  end

  // ===== Pipe stage 25:
  wire [31:0] p25_add_66407_comb;
  wire [31:0] p25_and_66450_comb;
  wire [31:0] p25_add_66429_comb;
  wire [31:0] p25_add_66431_comb;
  wire [31:0] p25_add_66454_comb;
  wire [31:0] p25_add_66432_comb;
  wire [31:0] p25_add_66433_comb;
  wire [31:0] p25_add_66455_comb;
  assign p25_add_66407_comb = p24_add_65894 + p24_add_66333;
  assign p25_and_66450_comb = p24_add_66356 & p24_add_66240;
  assign p25_add_66429_comb = {p25_add_66407_comb[5:0] ^ p25_add_66407_comb[10:5] ^ p25_add_66407_comb[24:19], p25_add_66407_comb[31:27] ^ p25_add_66407_comb[4:0] ^ p25_add_66407_comb[18:14], p25_add_66407_comb[26:13] ^ p25_add_66407_comb[31:18] ^ p25_add_66407_comb[13:0], p25_add_66407_comb[12:6] ^ p25_add_66407_comb[17:11] ^ p25_add_66407_comb[31:25]} + (p25_add_66407_comb & p24_add_66308 ^ ~(p25_add_66407_comb | ~p24_add_66192));
  assign p25_add_66431_comb = p25_add_66429_comb + 32'hd5a7_9147;
  assign p25_add_66454_comb = {p24_add_66356[1:0] ^ p24_add_66356[12:11] ^ p24_add_66356[21:20], p24_add_66356[31:21] ^ p24_add_66356[10:0] ^ p24_add_66356[19:9], p24_add_66356[20:12] ^ p24_add_66356[31:23] ^ p24_add_66356[8:0], p24_add_66356[11:2] ^ p24_add_66356[22:13] ^ p24_add_66356[31:22]} + (p25_and_66450_comb ^ p24_add_66356 & p24_add_66089 ^ p24_and_66351);
  assign p25_add_66432_comb = p25_add_66431_comb + p24_add_66334;
  assign p25_add_66433_comb = p24_add_66192 + p24_add_65690;
  assign p25_add_66455_comb = p24_add_66333 + p25_add_66454_comb;

  // Registers for pipe stage 25:
  reg [31:0] p25_add_66308;
  reg [31:0] p25_add_66407;
  reg [31:0] p25_add_66089;
  reg [31:0] p25_add_66432;
  reg [31:0] p25_add_66433;
  reg [31:0] p25_add_66240;
  reg [31:0] p25_add_66356;
  reg [31:0] p25_and_66450;
  reg [31:0] p25_add_66455;
  reg [31:0] p25_add_66257;
  reg [31:0] p25_add_66141;
  reg [31:0] p25_add_66124;
  reg [31:0] p25_add_66118;
  reg [31:0] p25_add_65794;
  reg [31:0] p25_add_65966;
  reg [31:0] p25_add_65760;
  reg [31:0] p25_add_65948;
  reg [31:0] p25_add_65524;
  reg [31:0] p25_add_65726;
  reg [31:0] p25_add_65930;
  reg [31:0] p25_add_65708;
  reg [31:0] p25_add_65912;
  reg [31:0] p25_add_65456;
  reg [31:0] p25_add_65690;
  reg [31:0] p25_add_64692;
  always_ff @ (posedge clk) begin
    p25_add_66308 <= p24_add_66308;
    p25_add_66407 <= p25_add_66407_comb;
    p25_add_66089 <= p24_add_66089;
    p25_add_66432 <= p25_add_66432_comb;
    p25_add_66433 <= p25_add_66433_comb;
    p25_add_66240 <= p24_add_66240;
    p25_add_66356 <= p24_add_66356;
    p25_and_66450 <= p25_and_66450_comb;
    p25_add_66455 <= p25_add_66455_comb;
    p25_add_66257 <= p24_add_66257;
    p25_add_66141 <= p24_add_66141;
    p25_add_66124 <= p24_add_66124;
    p25_add_66118 <= p24_add_66118;
    p25_add_65794 <= p24_add_65794;
    p25_add_65966 <= p24_add_65966;
    p25_add_65760 <= p24_add_65760;
    p25_add_65948 <= p24_add_65948;
    p25_add_65524 <= p24_add_65524;
    p25_add_65726 <= p24_add_65726;
    p25_add_65930 <= p24_add_65930;
    p25_add_65708 <= p24_add_65708;
    p25_add_65912 <= p24_add_65912;
    p25_add_65456 <= p24_add_65456;
    p25_add_65690 <= p24_add_65690;
    p25_add_64692 <= p24_add_64692;
  end

  // ===== Pipe stage 26:
  wire [31:0] p26_add_66506_comb;
  wire [31:0] p26_and_66549_comb;
  wire [31:0] p26_add_66528_comb;
  wire [31:0] p26_add_66530_comb;
  wire [31:0] p26_add_66553_comb;
  wire [31:0] p26_add_66531_comb;
  wire [31:0] p26_add_66532_comb;
  wire [31:0] p26_add_66554_comb;
  assign p26_add_66506_comb = p25_add_66089 + p25_add_66432;
  assign p26_and_66549_comb = p25_add_66455 & p25_add_66356;
  assign p26_add_66528_comb = {p26_add_66506_comb[5:0] ^ p26_add_66506_comb[10:5] ^ p26_add_66506_comb[24:19], p26_add_66506_comb[31:27] ^ p26_add_66506_comb[4:0] ^ p26_add_66506_comb[18:14], p26_add_66506_comb[26:13] ^ p26_add_66506_comb[31:18] ^ p26_add_66506_comb[13:0], p26_add_66506_comb[12:6] ^ p26_add_66506_comb[17:11] ^ p26_add_66506_comb[31:25]} + (p26_add_66506_comb & p25_add_66407 ^ ~(p26_add_66506_comb | ~p25_add_66308));
  assign p26_add_66530_comb = p26_add_66528_comb + 32'h06ca_6351;
  assign p26_add_66553_comb = {p25_add_66455[1:0] ^ p25_add_66455[12:11] ^ p25_add_66455[21:20], p25_add_66455[31:21] ^ p25_add_66455[10:0] ^ p25_add_66455[19:9], p25_add_66455[20:12] ^ p25_add_66455[31:23] ^ p25_add_66455[8:0], p25_add_66455[11:2] ^ p25_add_66455[22:13] ^ p25_add_66455[31:22]} + (p26_and_66549_comb ^ p25_add_66455 & p25_add_66240 ^ p25_and_66450);
  assign p26_add_66531_comb = p26_add_66530_comb + p25_add_66433;
  assign p26_add_66532_comb = p25_add_66308 + p25_add_65456;
  assign p26_add_66554_comb = p25_add_66432 + p26_add_66553_comb;

  // Registers for pipe stage 26:
  reg [31:0] p26_add_66407;
  reg [31:0] p26_add_66506;
  reg [31:0] p26_add_66240;
  reg [31:0] p26_add_66531;
  reg [31:0] p26_add_66532;
  reg [31:0] p26_add_66356;
  reg [31:0] p26_add_66455;
  reg [31:0] p26_and_66549;
  reg [31:0] p26_add_66554;
  reg [31:0] p26_add_66257;
  reg [31:0] p26_add_66141;
  reg [31:0] p26_add_66124;
  reg [31:0] p26_add_66118;
  reg [31:0] p26_add_65794;
  reg [31:0] p26_add_65966;
  reg [31:0] p26_add_65760;
  reg [31:0] p26_add_65948;
  reg [31:0] p26_add_65524;
  reg [31:0] p26_add_65726;
  reg [31:0] p26_add_65930;
  reg [31:0] p26_add_65708;
  reg [31:0] p26_add_65912;
  reg [31:0] p26_add_65456;
  reg [31:0] p26_add_65690;
  reg [31:0] p26_add_64692;
  always_ff @ (posedge clk) begin
    p26_add_66407 <= p25_add_66407;
    p26_add_66506 <= p26_add_66506_comb;
    p26_add_66240 <= p25_add_66240;
    p26_add_66531 <= p26_add_66531_comb;
    p26_add_66532 <= p26_add_66532_comb;
    p26_add_66356 <= p25_add_66356;
    p26_add_66455 <= p25_add_66455;
    p26_and_66549 <= p26_and_66549_comb;
    p26_add_66554 <= p26_add_66554_comb;
    p26_add_66257 <= p25_add_66257;
    p26_add_66141 <= p25_add_66141;
    p26_add_66124 <= p25_add_66124;
    p26_add_66118 <= p25_add_66118;
    p26_add_65794 <= p25_add_65794;
    p26_add_65966 <= p25_add_65966;
    p26_add_65760 <= p25_add_65760;
    p26_add_65948 <= p25_add_65948;
    p26_add_65524 <= p25_add_65524;
    p26_add_65726 <= p25_add_65726;
    p26_add_65930 <= p25_add_65930;
    p26_add_65708 <= p25_add_65708;
    p26_add_65912 <= p25_add_65912;
    p26_add_65456 <= p25_add_65456;
    p26_add_65690 <= p25_add_65690;
    p26_add_64692 <= p25_add_64692;
  end

  // ===== Pipe stage 27:
  wire [31:0] p27_add_66605_comb;
  wire [31:0] p27_and_66648_comb;
  wire [31:0] p27_add_66627_comb;
  wire [31:0] p27_add_66629_comb;
  wire [31:0] p27_add_66652_comb;
  wire [31:0] p27_add_66630_comb;
  wire [31:0] p27_add_66631_comb;
  wire [31:0] p27_add_66653_comb;
  assign p27_add_66605_comb = p26_add_66240 + p26_add_66531;
  assign p27_and_66648_comb = p26_add_66554 & p26_add_66455;
  assign p27_add_66627_comb = {p27_add_66605_comb[5:0] ^ p27_add_66605_comb[10:5] ^ p27_add_66605_comb[24:19], p27_add_66605_comb[31:27] ^ p27_add_66605_comb[4:0] ^ p27_add_66605_comb[18:14], p27_add_66605_comb[26:13] ^ p27_add_66605_comb[31:18] ^ p27_add_66605_comb[13:0], p27_add_66605_comb[12:6] ^ p27_add_66605_comb[17:11] ^ p27_add_66605_comb[31:25]} + (p27_add_66605_comb & p26_add_66506 ^ ~(p27_add_66605_comb | ~p26_add_66407));
  assign p27_add_66629_comb = p27_add_66627_comb + 32'h1429_2967;
  assign p27_add_66652_comb = {p26_add_66554[1:0] ^ p26_add_66554[12:11] ^ p26_add_66554[21:20], p26_add_66554[31:21] ^ p26_add_66554[10:0] ^ p26_add_66554[19:9], p26_add_66554[20:12] ^ p26_add_66554[31:23] ^ p26_add_66554[8:0], p26_add_66554[11:2] ^ p26_add_66554[22:13] ^ p26_add_66554[31:22]} + (p27_and_66648_comb ^ p26_add_66554 & p26_add_66356 ^ p26_and_66549);
  assign p27_add_66630_comb = p27_add_66629_comb + p26_add_66532;
  assign p27_add_66631_comb = p26_add_66407 + p26_add_65912;
  assign p27_add_66653_comb = p26_add_66531 + p27_add_66652_comb;

  // Registers for pipe stage 27:
  reg [31:0] p27_add_66506;
  reg [31:0] p27_add_66605;
  reg [31:0] p27_add_66356;
  reg [31:0] p27_add_66630;
  reg [31:0] p27_add_66631;
  reg [31:0] p27_add_66455;
  reg [31:0] p27_add_66554;
  reg [31:0] p27_and_66648;
  reg [31:0] p27_add_66653;
  reg [31:0] p27_add_66257;
  reg [31:0] p27_add_66141;
  reg [31:0] p27_add_66124;
  reg [31:0] p27_add_66118;
  reg [31:0] p27_add_65794;
  reg [31:0] p27_add_65966;
  reg [31:0] p27_add_65760;
  reg [31:0] p27_add_65948;
  reg [31:0] p27_add_65524;
  reg [31:0] p27_add_65726;
  reg [31:0] p27_add_65930;
  reg [31:0] p27_add_65708;
  reg [31:0] p27_add_65912;
  reg [31:0] p27_add_65456;
  reg [31:0] p27_add_65690;
  reg [31:0] p27_add_64692;
  always_ff @ (posedge clk) begin
    p27_add_66506 <= p26_add_66506;
    p27_add_66605 <= p27_add_66605_comb;
    p27_add_66356 <= p26_add_66356;
    p27_add_66630 <= p27_add_66630_comb;
    p27_add_66631 <= p27_add_66631_comb;
    p27_add_66455 <= p26_add_66455;
    p27_add_66554 <= p26_add_66554;
    p27_and_66648 <= p27_and_66648_comb;
    p27_add_66653 <= p27_add_66653_comb;
    p27_add_66257 <= p26_add_66257;
    p27_add_66141 <= p26_add_66141;
    p27_add_66124 <= p26_add_66124;
    p27_add_66118 <= p26_add_66118;
    p27_add_65794 <= p26_add_65794;
    p27_add_65966 <= p26_add_65966;
    p27_add_65760 <= p26_add_65760;
    p27_add_65948 <= p26_add_65948;
    p27_add_65524 <= p26_add_65524;
    p27_add_65726 <= p26_add_65726;
    p27_add_65930 <= p26_add_65930;
    p27_add_65708 <= p26_add_65708;
    p27_add_65912 <= p26_add_65912;
    p27_add_65456 <= p26_add_65456;
    p27_add_65690 <= p26_add_65690;
    p27_add_64692 <= p26_add_64692;
  end

  // ===== Pipe stage 28:
  wire [31:0] p28_add_66704_comb;
  wire [31:0] p28_and_66746_comb;
  wire [31:0] p28_add_66726_comb;
  wire [31:0] p28_add_66728_comb;
  wire [31:0] p28_add_66750_comb;
  wire [31:0] p28_add_66729_comb;
  wire [31:0] p28_add_66751_comb;
  assign p28_add_66704_comb = p27_add_66356 + p27_add_66630;
  assign p28_and_66746_comb = p27_add_66653 & p27_add_66554;
  assign p28_add_66726_comb = {p28_add_66704_comb[5:0] ^ p28_add_66704_comb[10:5] ^ p28_add_66704_comb[24:19], p28_add_66704_comb[31:27] ^ p28_add_66704_comb[4:0] ^ p28_add_66704_comb[18:14], p28_add_66704_comb[26:13] ^ p28_add_66704_comb[31:18] ^ p28_add_66704_comb[13:0], p28_add_66704_comb[12:6] ^ p28_add_66704_comb[17:11] ^ p28_add_66704_comb[31:25]} + (p28_add_66704_comb & p27_add_66605 ^ ~(p28_add_66704_comb | ~p27_add_66506));
  assign p28_add_66728_comb = p28_add_66726_comb + 32'h27b7_0a85;
  assign p28_add_66750_comb = {p27_add_66653[1:0] ^ p27_add_66653[12:11] ^ p27_add_66653[21:20], p27_add_66653[31:21] ^ p27_add_66653[10:0] ^ p27_add_66653[19:9], p27_add_66653[20:12] ^ p27_add_66653[31:23] ^ p27_add_66653[8:0], p27_add_66653[11:2] ^ p27_add_66653[22:13] ^ p27_add_66653[31:22]} + (p28_and_66746_comb ^ p27_add_66653 & p27_add_66455 ^ p27_and_66648);
  assign p28_add_66729_comb = p28_add_66728_comb + p27_add_66631;
  assign p28_add_66751_comb = p27_add_66630 + p28_add_66750_comb;

  // Registers for pipe stage 28:
  reg [31:0] p28_add_66506;
  reg [31:0] p28_add_66605;
  reg [31:0] p28_add_66704;
  reg [31:0] p28_add_66455;
  reg [31:0] p28_add_66729;
  reg [31:0] p28_add_66554;
  reg [31:0] p28_add_66653;
  reg [31:0] p28_and_66746;
  reg [31:0] p28_add_66751;
  reg [31:0] p28_add_66257;
  reg [31:0] p28_add_66141;
  reg [31:0] p28_add_66124;
  reg [31:0] p28_add_66118;
  reg [31:0] p28_add_65794;
  reg [31:0] p28_add_65966;
  reg [31:0] p28_add_65760;
  reg [31:0] p28_add_65948;
  reg [31:0] p28_add_65524;
  reg [31:0] p28_add_65726;
  reg [31:0] p28_add_65930;
  reg [31:0] p28_add_65708;
  reg [31:0] p28_add_65912;
  reg [31:0] p28_add_65456;
  reg [31:0] p28_add_65690;
  reg [31:0] p28_add_64692;
  always_ff @ (posedge clk) begin
    p28_add_66506 <= p27_add_66506;
    p28_add_66605 <= p27_add_66605;
    p28_add_66704 <= p28_add_66704_comb;
    p28_add_66455 <= p27_add_66455;
    p28_add_66729 <= p28_add_66729_comb;
    p28_add_66554 <= p27_add_66554;
    p28_add_66653 <= p27_add_66653;
    p28_and_66746 <= p28_and_66746_comb;
    p28_add_66751 <= p28_add_66751_comb;
    p28_add_66257 <= p27_add_66257;
    p28_add_66141 <= p27_add_66141;
    p28_add_66124 <= p27_add_66124;
    p28_add_66118 <= p27_add_66118;
    p28_add_65794 <= p27_add_65794;
    p28_add_65966 <= p27_add_65966;
    p28_add_65760 <= p27_add_65760;
    p28_add_65948 <= p27_add_65948;
    p28_add_65524 <= p27_add_65524;
    p28_add_65726 <= p27_add_65726;
    p28_add_65930 <= p27_add_65930;
    p28_add_65708 <= p27_add_65708;
    p28_add_65912 <= p27_add_65912;
    p28_add_65456 <= p27_add_65456;
    p28_add_65690 <= p27_add_65690;
    p28_add_64692 <= p27_add_64692;
  end

  // ===== Pipe stage 29:
  wire [31:0] p29_and_66852_comb;
  wire [31:0] p29_add_66802_comb;
  wire [31:0] p29_add_66856_comb;
  wire [31:0] p29_add_66857_comb;
  wire [28:0] p29_add_66824_comb;
  wire [31:0] p29_and_66874_comb;
  wire [31:0] p29_add_66829_comb;
  wire [31:0] p29_add_66830_comb;
  wire [31:0] p29_add_66831_comb;
  wire [31:0] p29_add_66878_comb;
  wire [31:0] p29_add_66832_comb;
  wire [29:0] p29_add_66835_comb;
  wire [31:0] p29_add_66879_comb;
  assign p29_and_66852_comb = p28_add_66751 & p28_add_66653;
  assign p29_add_66802_comb = p28_add_66455 + p28_add_66729;
  assign p29_add_66856_comb = {p28_add_66751[1:0] ^ p28_add_66751[12:11] ^ p28_add_66751[21:20], p28_add_66751[31:21] ^ p28_add_66751[10:0] ^ p28_add_66751[19:9], p28_add_66751[20:12] ^ p28_add_66751[31:23] ^ p28_add_66751[8:0], p28_add_66751[11:2] ^ p28_add_66751[22:13] ^ p28_add_66751[31:22]} + (p29_and_66852_comb ^ p28_add_66751 & p28_add_66554 ^ p28_and_66746);
  assign p29_add_66857_comb = p28_add_66729 + p29_add_66856_comb;
  assign p29_add_66824_comb = p28_add_65708[31:3] + 29'h05c3_6427;
  assign p29_and_66874_comb = p29_add_66857_comb & p28_add_66751;
  assign p29_add_66829_comb = {p29_add_66802_comb[5:0] ^ p29_add_66802_comb[10:5] ^ p29_add_66802_comb[24:19], p29_add_66802_comb[31:27] ^ p29_add_66802_comb[4:0] ^ p29_add_66802_comb[18:14], p29_add_66802_comb[26:13] ^ p29_add_66802_comb[31:18] ^ p29_add_66802_comb[13:0], p29_add_66802_comb[12:6] ^ p29_add_66802_comb[17:11] ^ p29_add_66802_comb[31:25]} + p28_add_66506;
  assign p29_add_66830_comb = (p29_add_66802_comb & p28_add_66704 ^ ~(p29_add_66802_comb | ~p28_add_66605)) + {p29_add_66824_comb, p28_add_65708[2:0]};
  assign p29_add_66831_comb = p29_add_66829_comb + p29_add_66830_comb;
  assign p29_add_66878_comb = {p29_add_66857_comb[1:0] ^ p29_add_66857_comb[12:11] ^ p29_add_66857_comb[21:20], p29_add_66857_comb[31:21] ^ p29_add_66857_comb[10:0] ^ p29_add_66857_comb[19:9], p29_add_66857_comb[20:12] ^ p29_add_66857_comb[31:23] ^ p29_add_66857_comb[8:0], p29_add_66857_comb[11:2] ^ p29_add_66857_comb[22:13] ^ p29_add_66857_comb[31:22]} + (p29_and_66874_comb ^ p29_add_66857_comb & p28_add_66653 ^ p29_and_66852_comb);
  assign p29_add_66832_comb = p28_add_66554 + p29_add_66831_comb;
  assign p29_add_66835_comb = p28_add_65930[31:2] + 30'h134b_1b7f;
  assign p29_add_66879_comb = p29_add_66831_comb + p29_add_66878_comb;

  // Registers for pipe stage 29:
  reg [31:0] p29_add_66605;
  reg [31:0] p29_add_66704;
  reg [31:0] p29_add_66802;
  reg [31:0] p29_add_66832;
  reg [29:0] p29_add_66835;
  reg [31:0] p29_add_66653;
  reg [31:0] p29_add_66751;
  reg [31:0] p29_add_66857;
  reg [31:0] p29_and_66874;
  reg [31:0] p29_add_66879;
  reg [31:0] p29_add_66257;
  reg [31:0] p29_add_66141;
  reg [31:0] p29_add_66124;
  reg [31:0] p29_add_66118;
  reg [31:0] p29_add_65794;
  reg [31:0] p29_add_65966;
  reg [31:0] p29_add_65760;
  reg [31:0] p29_add_65948;
  reg [31:0] p29_add_65524;
  reg [31:0] p29_add_65726;
  reg [31:0] p29_add_65930;
  reg [31:0] p29_add_65708;
  reg [31:0] p29_add_65912;
  reg [31:0] p29_add_65456;
  reg [31:0] p29_add_65690;
  reg [31:0] p29_add_64692;
  always_ff @ (posedge clk) begin
    p29_add_66605 <= p28_add_66605;
    p29_add_66704 <= p28_add_66704;
    p29_add_66802 <= p29_add_66802_comb;
    p29_add_66832 <= p29_add_66832_comb;
    p29_add_66835 <= p29_add_66835_comb;
    p29_add_66653 <= p28_add_66653;
    p29_add_66751 <= p28_add_66751;
    p29_add_66857 <= p29_add_66857_comb;
    p29_and_66874 <= p29_and_66874_comb;
    p29_add_66879 <= p29_add_66879_comb;
    p29_add_66257 <= p28_add_66257;
    p29_add_66141 <= p28_add_66141;
    p29_add_66124 <= p28_add_66124;
    p29_add_66118 <= p28_add_66118;
    p29_add_65794 <= p28_add_65794;
    p29_add_65966 <= p28_add_65966;
    p29_add_65760 <= p28_add_65760;
    p29_add_65948 <= p28_add_65948;
    p29_add_65524 <= p28_add_65524;
    p29_add_65726 <= p28_add_65726;
    p29_add_65930 <= p28_add_65930;
    p29_add_65708 <= p28_add_65708;
    p29_add_65912 <= p28_add_65912;
    p29_add_65456 <= p28_add_65456;
    p29_add_65690 <= p28_add_65690;
    p29_add_64692 <= p28_add_64692;
  end

  // ===== Pipe stage 30:
  wire [31:0] p30_add_66955_comb;
  wire [31:0] p30_add_66956_comb;
  wire [31:0] p30_add_66957_comb;
  wire [31:0] p30_add_66958_comb;
  wire [31:0] p30_and_67015_comb;
  wire [31:0] p30_add_66997_comb;
  wire [31:0] p30_add_66998_comb;
  wire [31:0] p30_add_67019_comb;
  wire [31:0] p30_add_67037_comb;
  wire [31:0] p30_add_66990_comb;
  wire [31:0] p30_add_66995_comb;
  wire [31:0] p30_add_67020_comb;
  wire [31:0] p30_add_67072_comb;
  wire [31:0] p30_add_67055_comb;
  wire [31:0] p30_add_67038_comb;
  assign p30_add_66955_comb = {p29_add_66832[5:0] ^ p29_add_66832[10:5] ^ p29_add_66832[24:19], p29_add_66832[31:27] ^ p29_add_66832[4:0] ^ p29_add_66832[18:14], p29_add_66832[26:13] ^ p29_add_66832[31:18] ^ p29_add_66832[13:0], p29_add_66832[12:6] ^ p29_add_66832[17:11] ^ p29_add_66832[31:25]} + p29_add_66605;
  assign p30_add_66956_comb = (p29_add_66832 & p29_add_66802 ^ ~(p29_add_66832 | ~p29_add_66704)) + {p29_add_66835, p29_add_65930[1:0]};
  assign p30_add_66957_comb = p30_add_66955_comb + p30_add_66956_comb;
  assign p30_add_66958_comb = p29_add_66653 + p30_add_66957_comb;
  assign p30_and_67015_comb = p29_add_66879 & p29_add_66857;
  assign p30_add_66997_comb = p29_add_64692 + {p29_add_65930[16:7] ^ p29_add_65930[18:9], p29_add_65930[6:0] ^ p29_add_65930[8:2] ^ p29_add_65930[31:25], p29_add_65930[31:30] ^ p29_add_65930[1:0] ^ p29_add_65930[24:23], p29_add_65930[29:17] ^ p29_add_65930[31:19] ^ p29_add_65930[22:10]};
  assign p30_add_66998_comb = p29_add_65524 + p30_add_66997_comb;
  assign p30_add_67019_comb = {p29_add_66879[1:0] ^ p29_add_66879[12:11] ^ p29_add_66879[21:20], p29_add_66879[31:21] ^ p29_add_66879[10:0] ^ p29_add_66879[19:9], p29_add_66879[20:12] ^ p29_add_66879[31:23] ^ p29_add_66879[8:0], p29_add_66879[11:2] ^ p29_add_66879[22:13] ^ p29_add_66879[31:22]} + (p30_and_67015_comb ^ p29_add_66879 & p29_add_66751 ^ p29_and_66874);
  assign p30_add_67037_comb = p30_add_66998_comb + {p29_add_66118[16:7] ^ p29_add_66118[18:9], p29_add_66118[6:0] ^ p29_add_66118[8:2] ^ p29_add_66118[31:25], p29_add_66118[31:30] ^ p29_add_66118[1:0] ^ p29_add_66118[24:23], p29_add_66118[29:17] ^ p29_add_66118[31:19] ^ p29_add_66118[22:10]};
  assign p30_add_66990_comb = {p30_add_66958_comb[5:0] ^ p30_add_66958_comb[10:5] ^ p30_add_66958_comb[24:19], p30_add_66958_comb[31:27] ^ p30_add_66958_comb[4:0] ^ p30_add_66958_comb[18:14], p30_add_66958_comb[26:13] ^ p30_add_66958_comb[31:18] ^ p30_add_66958_comb[13:0], p30_add_66958_comb[12:6] ^ p30_add_66958_comb[17:11] ^ p30_add_66958_comb[31:25]} + (p30_add_66958_comb & p29_add_66832 ^ ~(p30_add_66958_comb | ~p29_add_66802));
  assign p30_add_66995_comb = p29_add_66704 + p29_add_65726;
  assign p30_add_67020_comb = p30_add_66957_comb + p30_add_67019_comb;
  assign p30_add_67072_comb = {p29_add_65456[6:4] ^ p29_add_65456[17:15], p29_add_65456[3:0] ^ p29_add_65456[14:11] ^ p29_add_65456[31:28], p29_add_65456[31:21] ^ p29_add_65456[10:0] ^ p29_add_65456[27:17], p29_add_65456[20:7] ^ p29_add_65456[31:18] ^ p29_add_65456[16:3]} + p29_add_65690;
  assign p30_add_67055_comb = {p29_add_65690[6:4] ^ p29_add_65690[17:15], p29_add_65690[3:0] ^ p29_add_65690[14:11] ^ p29_add_65690[31:28], p29_add_65690[31:21] ^ p29_add_65690[10:0] ^ p29_add_65690[27:17], p29_add_65690[20:7] ^ p29_add_65690[31:18] ^ p29_add_65690[16:3]} + p29_add_64692;
  assign p30_add_67038_comb = p29_add_66141 + p30_add_67037_comb;

  // Registers for pipe stage 30:
  reg [31:0] p30_add_66802;
  reg [31:0] p30_add_66832;
  reg [31:0] p30_add_66958;
  reg [31:0] p30_add_66990;
  reg [31:0] p30_add_66995;
  reg [31:0] p30_add_66751;
  reg [31:0] p30_add_66857;
  reg [31:0] p30_add_66879;
  reg [31:0] p30_and_67015;
  reg [31:0] p30_add_67020;
  reg [31:0] p30_add_67072;
  reg [31:0] p30_add_67055;
  reg [31:0] p30_add_66257;
  reg [31:0] p30_add_67038;
  reg [31:0] p30_add_66124;
  reg [31:0] p30_add_66118;
  reg [31:0] p30_add_65794;
  reg [31:0] p30_add_65966;
  reg [31:0] p30_add_65760;
  reg [31:0] p30_add_65948;
  reg [31:0] p30_add_66998;
  reg [31:0] p30_add_65726;
  reg [31:0] p30_add_65930;
  reg [31:0] p30_add_65708;
  reg [31:0] p30_add_65912;
  reg [31:0] p30_add_65456;
  always_ff @ (posedge clk) begin
    p30_add_66802 <= p29_add_66802;
    p30_add_66832 <= p29_add_66832;
    p30_add_66958 <= p30_add_66958_comb;
    p30_add_66990 <= p30_add_66990_comb;
    p30_add_66995 <= p30_add_66995_comb;
    p30_add_66751 <= p29_add_66751;
    p30_add_66857 <= p29_add_66857;
    p30_add_66879 <= p29_add_66879;
    p30_and_67015 <= p30_and_67015_comb;
    p30_add_67020 <= p30_add_67020_comb;
    p30_add_67072 <= p30_add_67072_comb;
    p30_add_67055 <= p30_add_67055_comb;
    p30_add_66257 <= p29_add_66257;
    p30_add_67038 <= p30_add_67038_comb;
    p30_add_66124 <= p29_add_66124;
    p30_add_66118 <= p29_add_66118;
    p30_add_65794 <= p29_add_65794;
    p30_add_65966 <= p29_add_65966;
    p30_add_65760 <= p29_add_65760;
    p30_add_65948 <= p29_add_65948;
    p30_add_66998 <= p30_add_66998_comb;
    p30_add_65726 <= p29_add_65726;
    p30_add_65930 <= p29_add_65930;
    p30_add_65708 <= p29_add_65708;
    p30_add_65912 <= p29_add_65912;
    p30_add_65456 <= p29_add_65456;
  end

  // ===== Pipe stage 31:
  wire [31:0] p31_add_67173_comb;
  wire [31:0] p31_add_67126_comb;
  wire [31:0] p31_add_67174_comb;
  wire [31:0] p31_add_67127_comb;
  wire [31:0] p31_add_67128_comb;
  wire [31:0] p31_and_67191_comb;
  wire [29:0] p31_add_67150_comb;
  wire [31:0] p31_add_67195_comb;
  wire [31:0] p31_add_67231_comb;
  wire [31:0] p31_add_67213_comb;
  wire [31:0] p31_add_67171_comb;
  wire [31:0] p31_add_67196_comb;
  wire [31:0] p31_add_67300_comb;
  wire [31:0] p31_add_67283_comb;
  wire [31:0] p31_add_67266_comb;
  wire [31:0] p31_add_67249_comb;
  wire [31:0] p31_add_67232_comb;
  wire [31:0] p31_add_67214_comb;
  wire [31:0] p31_add_67155_comb;
  wire [31:0] p31_add_67156_comb;
  assign p31_add_67173_comb = p30_add_65456 + {p30_add_66998[16:7] ^ p30_add_66998[18:9], p30_add_66998[6:0] ^ p30_add_66998[8:2] ^ p30_add_66998[31:25], p30_add_66998[31:30] ^ p30_add_66998[1:0] ^ p30_add_66998[24:23], p30_add_66998[29:17] ^ p30_add_66998[31:19] ^ p30_add_66998[22:10]};
  assign p31_add_67126_comb = p30_add_66990 + 32'h5338_0d13;
  assign p31_add_67174_comb = p30_add_65760 + p31_add_67173_comb;
  assign p31_add_67127_comb = p31_add_67126_comb + p30_add_66995;
  assign p31_add_67128_comb = p30_add_66751 + p31_add_67127_comb;
  assign p31_and_67191_comb = p30_add_67020 & p30_add_66879;
  assign p31_add_67150_comb = p30_add_66998[31:2] + 30'h1942_9cd5;
  assign p31_add_67195_comb = {p30_add_67020[1:0] ^ p30_add_67020[12:11] ^ p30_add_67020[21:20], p30_add_67020[31:21] ^ p30_add_67020[10:0] ^ p30_add_67020[19:9], p30_add_67020[20:12] ^ p30_add_67020[31:23] ^ p30_add_67020[8:0], p30_add_67020[11:2] ^ p30_add_67020[22:13] ^ p30_add_67020[31:22]} + (p31_and_67191_comb ^ p30_add_67020 & p30_add_66857 ^ p30_and_67015);
  assign p31_add_67231_comb = p31_add_67174_comb + {p30_add_67038[16:7] ^ p30_add_67038[18:9], p30_add_67038[6:0] ^ p30_add_67038[8:2] ^ p30_add_67038[31:25], p30_add_67038[31:30] ^ p30_add_67038[1:0] ^ p30_add_67038[24:23], p30_add_67038[29:17] ^ p30_add_67038[31:19] ^ p30_add_67038[22:10]};
  assign p31_add_67213_comb = p30_add_65708 + {p31_add_67174_comb[16:7] ^ p31_add_67174_comb[18:9], p31_add_67174_comb[6:0] ^ p31_add_67174_comb[8:2] ^ p31_add_67174_comb[31:25], p31_add_67174_comb[31:30] ^ p31_add_67174_comb[1:0] ^ p31_add_67174_comb[24:23], p31_add_67174_comb[29:17] ^ p31_add_67174_comb[31:19] ^ p31_add_67174_comb[22:10]};
  assign p31_add_67171_comb = p30_add_66832 + p30_add_65948;
  assign p31_add_67196_comb = p31_add_67127_comb + p31_add_67195_comb;
  assign p31_add_67300_comb = {p30_add_65726[6:4] ^ p30_add_65726[17:15], p30_add_65726[3:0] ^ p30_add_65726[14:11] ^ p30_add_65726[31:28], p30_add_65726[31:21] ^ p30_add_65726[10:0] ^ p30_add_65726[27:17], p30_add_65726[20:7] ^ p30_add_65726[31:18] ^ p30_add_65726[16:3]} + p30_add_65930;
  assign p31_add_67283_comb = {p30_add_65930[6:4] ^ p30_add_65930[17:15], p30_add_65930[3:0] ^ p30_add_65930[14:11] ^ p30_add_65930[31:28], p30_add_65930[31:21] ^ p30_add_65930[10:0] ^ p30_add_65930[27:17], p30_add_65930[20:7] ^ p30_add_65930[31:18] ^ p30_add_65930[16:3]} + p30_add_65708;
  assign p31_add_67266_comb = {p30_add_65708[6:4] ^ p30_add_65708[17:15], p30_add_65708[3:0] ^ p30_add_65708[14:11] ^ p30_add_65708[31:28], p30_add_65708[31:21] ^ p30_add_65708[10:0] ^ p30_add_65708[27:17], p30_add_65708[20:7] ^ p30_add_65708[31:18] ^ p30_add_65708[16:3]} + p30_add_65912;
  assign p31_add_67249_comb = {p30_add_65912[6:4] ^ p30_add_65912[17:15], p30_add_65912[3:0] ^ p30_add_65912[14:11] ^ p30_add_65912[31:28], p30_add_65912[31:21] ^ p30_add_65912[10:0] ^ p30_add_65912[27:17], p30_add_65912[20:7] ^ p30_add_65912[31:18] ^ p30_add_65912[16:3]} + p30_add_65456;
  assign p31_add_67232_comb = p30_add_67055 + p31_add_67231_comb;
  assign p31_add_67214_comb = p30_add_65794 + p31_add_67213_comb;
  assign p31_add_67155_comb = {p31_add_67128_comb[5:0] ^ p31_add_67128_comb[10:5] ^ p31_add_67128_comb[24:19], p31_add_67128_comb[31:27] ^ p31_add_67128_comb[4:0] ^ p31_add_67128_comb[18:14], p31_add_67128_comb[26:13] ^ p31_add_67128_comb[31:18] ^ p31_add_67128_comb[13:0], p31_add_67128_comb[12:6] ^ p31_add_67128_comb[17:11] ^ p31_add_67128_comb[31:25]} + p30_add_66802;
  assign p31_add_67156_comb = (p31_add_67128_comb & p30_add_66958 ^ ~(p31_add_67128_comb | ~p30_add_66832)) + {p31_add_67150_comb, p30_add_66998[1:0]};

  // Registers for pipe stage 31:
  reg [31:0] p31_add_66958;
  reg [31:0] p31_add_67128;
  reg [31:0] p31_add_66857;
  reg [31:0] p31_add_67171;
  reg [31:0] p31_add_66879;
  reg [31:0] p31_add_67020;
  reg [31:0] p31_and_67191;
  reg [31:0] p31_add_67196;
  reg [31:0] p31_add_67300;
  reg [31:0] p31_add_67283;
  reg [31:0] p31_add_67266;
  reg [31:0] p31_add_67249;
  reg [31:0] p31_add_67072;
  reg [31:0] p31_add_67232;
  reg [31:0] p31_add_66257;
  reg [31:0] p31_add_67038;
  reg [31:0] p31_add_66124;
  reg [31:0] p31_add_66118;
  reg [31:0] p31_add_67214;
  reg [31:0] p31_add_65966;
  reg [31:0] p31_add_67174;
  reg [31:0] p31_add_65948;
  reg [31:0] p31_add_67155;
  reg [31:0] p31_add_67156;
  reg [31:0] p31_add_66998;
  reg [31:0] p31_add_65726;
  always_ff @ (posedge clk) begin
    p31_add_66958 <= p30_add_66958;
    p31_add_67128 <= p31_add_67128_comb;
    p31_add_66857 <= p30_add_66857;
    p31_add_67171 <= p31_add_67171_comb;
    p31_add_66879 <= p30_add_66879;
    p31_add_67020 <= p30_add_67020;
    p31_and_67191 <= p31_and_67191_comb;
    p31_add_67196 <= p31_add_67196_comb;
    p31_add_67300 <= p31_add_67300_comb;
    p31_add_67283 <= p31_add_67283_comb;
    p31_add_67266 <= p31_add_67266_comb;
    p31_add_67249 <= p31_add_67249_comb;
    p31_add_67072 <= p30_add_67072;
    p31_add_67232 <= p31_add_67232_comb;
    p31_add_66257 <= p30_add_66257;
    p31_add_67038 <= p30_add_67038;
    p31_add_66124 <= p30_add_66124;
    p31_add_66118 <= p30_add_66118;
    p31_add_67214 <= p31_add_67214_comb;
    p31_add_65966 <= p30_add_65966;
    p31_add_67174 <= p31_add_67174_comb;
    p31_add_65948 <= p30_add_65948;
    p31_add_67155 <= p31_add_67155_comb;
    p31_add_67156 <= p31_add_67156_comb;
    p31_add_66998 <= p30_add_66998;
    p31_add_65726 <= p30_add_65726;
  end

  // ===== Pipe stage 32:
  wire [31:0] p32_add_67353_comb;
  wire [31:0] p32_add_67417_comb;
  wire [31:0] p32_add_67354_comb;
  wire [31:0] p32_add_67418_comb;
  wire [31:0] p32_and_67395_comb;
  wire [31:0] p32_add_67399_comb;
  wire [31:0] p32_add_67376_comb;
  wire [31:0] p32_add_67435_comb;
  wire [31:0] p32_add_67400_comb;
  wire [31:0] p32_add_67378_comb;
  wire [31:0] p32_add_67487_comb;
  wire [31:0] p32_add_67470_comb;
  wire [31:0] p32_add_67453_comb;
  wire [31:0] p32_add_67436_comb;
  assign p32_add_67353_comb = p31_add_67155 + p31_add_67156;
  assign p32_add_67417_comb = p31_add_65726 + {p31_add_67214[16:7] ^ p31_add_67214[18:9], p31_add_67214[6:0] ^ p31_add_67214[8:2] ^ p31_add_67214[31:25], p31_add_67214[31:30] ^ p31_add_67214[1:0] ^ p31_add_67214[24:23], p31_add_67214[29:17] ^ p31_add_67214[31:19] ^ p31_add_67214[22:10]};
  assign p32_add_67354_comb = p31_add_66857 + p32_add_67353_comb;
  assign p32_add_67418_comb = p31_add_66124 + p32_add_67417_comb;
  assign p32_and_67395_comb = p31_add_67196 & p31_add_67020;
  assign p32_add_67399_comb = {p31_add_67196[1:0] ^ p31_add_67196[12:11] ^ p31_add_67196[21:20], p31_add_67196[31:21] ^ p31_add_67196[10:0] ^ p31_add_67196[19:9], p31_add_67196[20:12] ^ p31_add_67196[31:23] ^ p31_add_67196[8:0], p31_add_67196[11:2] ^ p31_add_67196[22:13] ^ p31_add_67196[31:22]} + (p32_and_67395_comb ^ p31_add_67196 & p31_add_66879 ^ p31_and_67191);
  assign p32_add_67376_comb = {p32_add_67354_comb[5:0] ^ p32_add_67354_comb[10:5] ^ p32_add_67354_comb[24:19], p32_add_67354_comb[31:27] ^ p32_add_67354_comb[4:0] ^ p32_add_67354_comb[18:14], p32_add_67354_comb[26:13] ^ p32_add_67354_comb[31:18] ^ p32_add_67354_comb[13:0], p32_add_67354_comb[12:6] ^ p32_add_67354_comb[17:11] ^ p32_add_67354_comb[31:25]} + (p32_add_67354_comb & p31_add_67128 ^ ~(p32_add_67354_comb | ~p31_add_66958));
  assign p32_add_67435_comb = p31_add_65948 + {p32_add_67418_comb[16:7] ^ p32_add_67418_comb[18:9], p32_add_67418_comb[6:0] ^ p32_add_67418_comb[8:2] ^ p32_add_67418_comb[31:25], p32_add_67418_comb[31:30] ^ p32_add_67418_comb[1:0] ^ p32_add_67418_comb[24:23], p32_add_67418_comb[29:17] ^ p32_add_67418_comb[31:19] ^ p32_add_67418_comb[22:10]};
  assign p32_add_67400_comb = p32_add_67353_comb + p32_add_67399_comb;
  assign p32_add_67378_comb = p32_add_67376_comb + 32'h766a_0abb;
  assign p32_add_67487_comb = {p31_add_67174[6:4] ^ p31_add_67174[17:15], p31_add_67174[3:0] ^ p31_add_67174[14:11] ^ p31_add_67174[31:28], p31_add_67174[31:21] ^ p31_add_67174[10:0] ^ p31_add_67174[27:17], p31_add_67174[20:7] ^ p31_add_67174[31:18] ^ p31_add_67174[16:3]} + p31_add_65948;
  assign p32_add_67470_comb = {p31_add_65948[6:4] ^ p31_add_65948[17:15], p31_add_65948[3:0] ^ p31_add_65948[14:11] ^ p31_add_65948[31:28], p31_add_65948[31:21] ^ p31_add_65948[10:0] ^ p31_add_65948[27:17], p31_add_65948[20:7] ^ p31_add_65948[31:18] ^ p31_add_65948[16:3]} + p31_add_66998;
  assign p32_add_67453_comb = {p31_add_66998[6:4] ^ p31_add_66998[17:15], p31_add_66998[3:0] ^ p31_add_66998[14:11] ^ p31_add_66998[31:28], p31_add_66998[31:21] ^ p31_add_66998[10:0] ^ p31_add_66998[27:17], p31_add_66998[20:7] ^ p31_add_66998[31:18] ^ p31_add_66998[16:3]} + p31_add_65726;
  assign p32_add_67436_comb = p31_add_66257 + p32_add_67435_comb;

  // Registers for pipe stage 32:
  reg [31:0] p32_add_66958;
  reg [31:0] p32_add_67128;
  reg [31:0] p32_add_67354;
  reg [31:0] p32_add_67171;
  reg [31:0] p32_add_66879;
  reg [31:0] p32_add_67020;
  reg [31:0] p32_add_67196;
  reg [31:0] p32_and_67395;
  reg [31:0] p32_add_67400;
  reg [31:0] p32_add_67378;
  reg [31:0] p32_add_67487;
  reg [31:0] p32_add_67470;
  reg [31:0] p32_add_67453;
  reg [31:0] p32_add_67300;
  reg [31:0] p32_add_67283;
  reg [31:0] p32_add_67266;
  reg [31:0] p32_add_67249;
  reg [31:0] p32_add_67072;
  reg [31:0] p32_add_67232;
  reg [31:0] p32_add_67436;
  reg [31:0] p32_add_67038;
  reg [31:0] p32_add_67418;
  reg [31:0] p32_add_66118;
  reg [31:0] p32_add_67214;
  reg [31:0] p32_add_65966;
  reg [31:0] p32_add_67174;
  always_ff @ (posedge clk) begin
    p32_add_66958 <= p31_add_66958;
    p32_add_67128 <= p31_add_67128;
    p32_add_67354 <= p32_add_67354_comb;
    p32_add_67171 <= p31_add_67171;
    p32_add_66879 <= p31_add_66879;
    p32_add_67020 <= p31_add_67020;
    p32_add_67196 <= p31_add_67196;
    p32_and_67395 <= p32_and_67395_comb;
    p32_add_67400 <= p32_add_67400_comb;
    p32_add_67378 <= p32_add_67378_comb;
    p32_add_67487 <= p32_add_67487_comb;
    p32_add_67470 <= p32_add_67470_comb;
    p32_add_67453 <= p32_add_67453_comb;
    p32_add_67300 <= p31_add_67300;
    p32_add_67283 <= p31_add_67283;
    p32_add_67266 <= p31_add_67266;
    p32_add_67249 <= p31_add_67249;
    p32_add_67072 <= p31_add_67072;
    p32_add_67232 <= p31_add_67232;
    p32_add_67436 <= p32_add_67436_comb;
    p32_add_67038 <= p31_add_67038;
    p32_add_67418 <= p32_add_67418_comb;
    p32_add_66118 <= p31_add_66118;
    p32_add_67214 <= p31_add_67214;
    p32_add_65966 <= p31_add_65966;
    p32_add_67174 <= p31_add_67174;
  end

  // ===== Pipe stage 33:
  wire [31:0] p33_add_67610_comb;
  wire [31:0] p33_add_67540_comb;
  wire [31:0] p33_add_67611_comb;
  wire [31:0] p33_add_67541_comb;
  wire [31:0] p33_and_67588_comb;
  wire [30:0] p33_add_67563_comb;
  wire [31:0] p33_add_67592_comb;
  wire [31:0] p33_add_67628_comb;
  wire [31:0] p33_add_67568_comb;
  wire [31:0] p33_add_67569_comb;
  wire [31:0] p33_add_67571_comb;
  wire [31:0] p33_add_67593_comb;
  wire [31:0] p33_add_67663_comb;
  wire [31:0] p33_add_67646_comb;
  wire [31:0] p33_add_67629_comb;
  wire [31:0] p33_add_67570_comb;
  assign p33_add_67610_comb = p32_add_65966 + {p32_add_67436[16:7] ^ p32_add_67436[18:9], p32_add_67436[6:0] ^ p32_add_67436[8:2] ^ p32_add_67436[31:25], p32_add_67436[31:30] ^ p32_add_67436[1:0] ^ p32_add_67436[24:23], p32_add_67436[29:17] ^ p32_add_67436[31:19] ^ p32_add_67436[22:10]};
  assign p33_add_67540_comb = p32_add_67378 + p32_add_67171;
  assign p33_add_67611_comb = p32_add_67072 + p33_add_67610_comb;
  assign p33_add_67541_comb = p32_add_66879 + p33_add_67540_comb;
  assign p33_and_67588_comb = p32_add_67400 & p32_add_67196;
  assign p33_add_67563_comb = p32_add_67174[31:1] + 31'h40e1_6497;
  assign p33_add_67592_comb = {p32_add_67400[1:0] ^ p32_add_67400[12:11] ^ p32_add_67400[21:20], p32_add_67400[31:21] ^ p32_add_67400[10:0] ^ p32_add_67400[19:9], p32_add_67400[20:12] ^ p32_add_67400[31:23] ^ p32_add_67400[8:0], p32_add_67400[11:2] ^ p32_add_67400[22:13] ^ p32_add_67400[31:22]} + (p33_and_67588_comb ^ p32_add_67400 & p32_add_67020 ^ p32_and_67395);
  assign p33_add_67628_comb = p32_add_66118 + {p33_add_67611_comb[16:7] ^ p33_add_67611_comb[18:9], p33_add_67611_comb[6:0] ^ p33_add_67611_comb[8:2] ^ p33_add_67611_comb[31:25], p33_add_67611_comb[31:30] ^ p33_add_67611_comb[1:0] ^ p33_add_67611_comb[24:23], p33_add_67611_comb[29:17] ^ p33_add_67611_comb[31:19] ^ p33_add_67611_comb[22:10]};
  assign p33_add_67568_comb = {p33_add_67541_comb[5:0] ^ p33_add_67541_comb[10:5] ^ p33_add_67541_comb[24:19], p33_add_67541_comb[31:27] ^ p33_add_67541_comb[4:0] ^ p33_add_67541_comb[18:14], p33_add_67541_comb[26:13] ^ p33_add_67541_comb[31:18] ^ p33_add_67541_comb[13:0], p33_add_67541_comb[12:6] ^ p33_add_67541_comb[17:11] ^ p33_add_67541_comb[31:25]} + p32_add_66958;
  assign p33_add_67569_comb = (p33_add_67541_comb & p32_add_67354 ^ ~(p33_add_67541_comb | ~p32_add_67128)) + {p33_add_67563_comb, p32_add_67174[0]};
  assign p33_add_67571_comb = p32_add_67128 + p32_add_65966;
  assign p33_add_67593_comb = p33_add_67540_comb + p33_add_67592_comb;
  assign p33_add_67663_comb = {p32_add_67214[6:4] ^ p32_add_67214[17:15], p32_add_67214[3:0] ^ p32_add_67214[14:11] ^ p32_add_67214[31:28], p32_add_67214[31:21] ^ p32_add_67214[10:0] ^ p32_add_67214[27:17], p32_add_67214[20:7] ^ p32_add_67214[31:18] ^ p32_add_67214[16:3]} + p32_add_65966;
  assign p33_add_67646_comb = {p32_add_65966[6:4] ^ p32_add_65966[17:15], p32_add_65966[3:0] ^ p32_add_65966[14:11] ^ p32_add_65966[31:28], p32_add_65966[31:21] ^ p32_add_65966[10:0] ^ p32_add_65966[27:17], p32_add_65966[20:7] ^ p32_add_65966[31:18] ^ p32_add_65966[16:3]} + p32_add_67174;
  assign p33_add_67629_comb = p32_add_67266 + p33_add_67628_comb;
  assign p33_add_67570_comb = p33_add_67568_comb + p33_add_67569_comb;

  // Registers for pipe stage 33:
  reg [31:0] p33_add_67354;
  reg [31:0] p33_add_67541;
  reg [31:0] p33_add_67020;
  reg [31:0] p33_add_67571;
  reg [31:0] p33_add_67196;
  reg [31:0] p33_add_67400;
  reg [31:0] p33_and_67588;
  reg [31:0] p33_add_67593;
  reg [31:0] p33_add_67663;
  reg [31:0] p33_add_67646;
  reg [31:0] p33_add_67487;
  reg [31:0] p33_add_67470;
  reg [31:0] p33_add_67453;
  reg [31:0] p33_add_67300;
  reg [31:0] p33_add_67283;
  reg [31:0] p33_add_67629;
  reg [31:0] p33_add_67249;
  reg [31:0] p33_add_67611;
  reg [31:0] p33_add_67232;
  reg [31:0] p33_add_67436;
  reg [31:0] p33_add_67038;
  reg [31:0] p33_add_67418;
  reg [31:0] p33_add_66118;
  reg [31:0] p33_add_67214;
  reg [31:0] p33_add_67570;
  always_ff @ (posedge clk) begin
    p33_add_67354 <= p32_add_67354;
    p33_add_67541 <= p33_add_67541_comb;
    p33_add_67020 <= p32_add_67020;
    p33_add_67571 <= p33_add_67571_comb;
    p33_add_67196 <= p32_add_67196;
    p33_add_67400 <= p32_add_67400;
    p33_and_67588 <= p33_and_67588_comb;
    p33_add_67593 <= p33_add_67593_comb;
    p33_add_67663 <= p33_add_67663_comb;
    p33_add_67646 <= p33_add_67646_comb;
    p33_add_67487 <= p32_add_67487;
    p33_add_67470 <= p32_add_67470;
    p33_add_67453 <= p32_add_67453;
    p33_add_67300 <= p32_add_67300;
    p33_add_67283 <= p32_add_67283;
    p33_add_67629 <= p33_add_67629_comb;
    p33_add_67249 <= p32_add_67249;
    p33_add_67611 <= p33_add_67611_comb;
    p33_add_67232 <= p32_add_67232;
    p33_add_67436 <= p32_add_67436;
    p33_add_67038 <= p32_add_67038;
    p33_add_67418 <= p32_add_67418;
    p33_add_66118 <= p32_add_66118;
    p33_add_67214 <= p32_add_67214;
    p33_add_67570 <= p33_add_67570_comb;
  end

  // ===== Pipe stage 34:
  wire [31:0] p34_add_67714_comb;
  wire [31:0] p34_and_67757_comb;
  wire [31:0] p34_add_67736_comb;
  wire [31:0] p34_add_67738_comb;
  wire [31:0] p34_add_67761_comb;
  wire [31:0] p34_add_67779_comb;
  wire [31:0] p34_add_67739_comb;
  wire [31:0] p34_add_67740_comb;
  wire [31:0] p34_add_67762_comb;
  wire [31:0] p34_add_67780_comb;
  assign p34_add_67714_comb = p33_add_67020 + p33_add_67570;
  assign p34_and_67757_comb = p33_add_67593 & p33_add_67400;
  assign p34_add_67736_comb = {p34_add_67714_comb[5:0] ^ p34_add_67714_comb[10:5] ^ p34_add_67714_comb[24:19], p34_add_67714_comb[31:27] ^ p34_add_67714_comb[4:0] ^ p34_add_67714_comb[18:14], p34_add_67714_comb[26:13] ^ p34_add_67714_comb[31:18] ^ p34_add_67714_comb[13:0], p34_add_67714_comb[12:6] ^ p34_add_67714_comb[17:11] ^ p34_add_67714_comb[31:25]} + (p34_add_67714_comb & p33_add_67541 ^ ~(p34_add_67714_comb | ~p33_add_67354));
  assign p34_add_67738_comb = p34_add_67736_comb + 32'h9272_2c85;
  assign p34_add_67761_comb = {p33_add_67593[1:0] ^ p33_add_67593[12:11] ^ p33_add_67593[21:20], p33_add_67593[31:21] ^ p33_add_67593[10:0] ^ p33_add_67593[19:9], p33_add_67593[20:12] ^ p33_add_67593[31:23] ^ p33_add_67593[8:0], p33_add_67593[11:2] ^ p33_add_67593[22:13] ^ p33_add_67593[31:22]} + (p34_and_67757_comb ^ p33_add_67593 & p33_add_67196 ^ p33_and_67588);
  assign p34_add_67779_comb = p33_add_67038 + {p33_add_67629[16:7] ^ p33_add_67629[18:9], p33_add_67629[6:0] ^ p33_add_67629[8:2] ^ p33_add_67629[31:25], p33_add_67629[31:30] ^ p33_add_67629[1:0] ^ p33_add_67629[24:23], p33_add_67629[29:17] ^ p33_add_67629[31:19] ^ p33_add_67629[22:10]};
  assign p34_add_67739_comb = p34_add_67738_comb + p33_add_67571;
  assign p34_add_67740_comb = p33_add_67354 + p33_add_67214;
  assign p34_add_67762_comb = p33_add_67570 + p34_add_67761_comb;
  assign p34_add_67780_comb = p33_add_67300 + p34_add_67779_comb;

  // Registers for pipe stage 34:
  reg [31:0] p34_add_67541;
  reg [31:0] p34_add_67714;
  reg [31:0] p34_add_67196;
  reg [31:0] p34_add_67739;
  reg [31:0] p34_add_67740;
  reg [31:0] p34_add_67400;
  reg [31:0] p34_add_67593;
  reg [31:0] p34_and_67757;
  reg [31:0] p34_add_67762;
  reg [31:0] p34_add_67663;
  reg [31:0] p34_add_67646;
  reg [31:0] p34_add_67487;
  reg [31:0] p34_add_67470;
  reg [31:0] p34_add_67453;
  reg [31:0] p34_add_67780;
  reg [31:0] p34_add_67283;
  reg [31:0] p34_add_67629;
  reg [31:0] p34_add_67249;
  reg [31:0] p34_add_67611;
  reg [31:0] p34_add_67232;
  reg [31:0] p34_add_67436;
  reg [31:0] p34_add_67038;
  reg [31:0] p34_add_67418;
  reg [31:0] p34_add_66118;
  reg [31:0] p34_add_67214;
  always_ff @ (posedge clk) begin
    p34_add_67541 <= p33_add_67541;
    p34_add_67714 <= p34_add_67714_comb;
    p34_add_67196 <= p33_add_67196;
    p34_add_67739 <= p34_add_67739_comb;
    p34_add_67740 <= p34_add_67740_comb;
    p34_add_67400 <= p33_add_67400;
    p34_add_67593 <= p33_add_67593;
    p34_and_67757 <= p34_and_67757_comb;
    p34_add_67762 <= p34_add_67762_comb;
    p34_add_67663 <= p33_add_67663;
    p34_add_67646 <= p33_add_67646;
    p34_add_67487 <= p33_add_67487;
    p34_add_67470 <= p33_add_67470;
    p34_add_67453 <= p33_add_67453;
    p34_add_67780 <= p34_add_67780_comb;
    p34_add_67283 <= p33_add_67283;
    p34_add_67629 <= p33_add_67629;
    p34_add_67249 <= p33_add_67249;
    p34_add_67611 <= p33_add_67611;
    p34_add_67232 <= p33_add_67232;
    p34_add_67436 <= p33_add_67436;
    p34_add_67038 <= p33_add_67038;
    p34_add_67418 <= p33_add_67418;
    p34_add_66118 <= p33_add_66118;
    p34_add_67214 <= p33_add_67214;
  end

  // ===== Pipe stage 35:
  wire [31:0] p35_add_67831_comb;
  wire [31:0] p35_and_67874_comb;
  wire [31:0] p35_add_67853_comb;
  wire [31:0] p35_add_67855_comb;
  wire [31:0] p35_add_67878_comb;
  wire [31:0] p35_add_67856_comb;
  wire [31:0] p35_add_67857_comb;
  wire [31:0] p35_add_67879_comb;
  assign p35_add_67831_comb = p34_add_67196 + p34_add_67739;
  assign p35_and_67874_comb = p34_add_67762 & p34_add_67593;
  assign p35_add_67853_comb = {p35_add_67831_comb[5:0] ^ p35_add_67831_comb[10:5] ^ p35_add_67831_comb[24:19], p35_add_67831_comb[31:27] ^ p35_add_67831_comb[4:0] ^ p35_add_67831_comb[18:14], p35_add_67831_comb[26:13] ^ p35_add_67831_comb[31:18] ^ p35_add_67831_comb[13:0], p35_add_67831_comb[12:6] ^ p35_add_67831_comb[17:11] ^ p35_add_67831_comb[31:25]} + (p35_add_67831_comb & p34_add_67714 ^ ~(p35_add_67831_comb | ~p34_add_67541));
  assign p35_add_67855_comb = p35_add_67853_comb + 32'ha2bf_e8a1;
  assign p35_add_67878_comb = {p34_add_67762[1:0] ^ p34_add_67762[12:11] ^ p34_add_67762[21:20], p34_add_67762[31:21] ^ p34_add_67762[10:0] ^ p34_add_67762[19:9], p34_add_67762[20:12] ^ p34_add_67762[31:23] ^ p34_add_67762[8:0], p34_add_67762[11:2] ^ p34_add_67762[22:13] ^ p34_add_67762[31:22]} + (p35_and_67874_comb ^ p34_add_67762 & p34_add_67400 ^ p34_and_67757);
  assign p35_add_67856_comb = p35_add_67855_comb + p34_add_67740;
  assign p35_add_67857_comb = p34_add_67541 + p34_add_66118;
  assign p35_add_67879_comb = p34_add_67739 + p35_add_67878_comb;

  // Registers for pipe stage 35:
  reg [31:0] p35_add_67714;
  reg [31:0] p35_add_67831;
  reg [31:0] p35_add_67400;
  reg [31:0] p35_add_67856;
  reg [31:0] p35_add_67857;
  reg [31:0] p35_add_67593;
  reg [31:0] p35_add_67762;
  reg [31:0] p35_and_67874;
  reg [31:0] p35_add_67879;
  reg [31:0] p35_add_67663;
  reg [31:0] p35_add_67646;
  reg [31:0] p35_add_67487;
  reg [31:0] p35_add_67470;
  reg [31:0] p35_add_67453;
  reg [31:0] p35_add_67780;
  reg [31:0] p35_add_67283;
  reg [31:0] p35_add_67629;
  reg [31:0] p35_add_67249;
  reg [31:0] p35_add_67611;
  reg [31:0] p35_add_67232;
  reg [31:0] p35_add_67436;
  reg [31:0] p35_add_67038;
  reg [31:0] p35_add_67418;
  reg [31:0] p35_add_66118;
  reg [31:0] p35_add_67214;
  always_ff @ (posedge clk) begin
    p35_add_67714 <= p34_add_67714;
    p35_add_67831 <= p35_add_67831_comb;
    p35_add_67400 <= p34_add_67400;
    p35_add_67856 <= p35_add_67856_comb;
    p35_add_67857 <= p35_add_67857_comb;
    p35_add_67593 <= p34_add_67593;
    p35_add_67762 <= p34_add_67762;
    p35_and_67874 <= p35_and_67874_comb;
    p35_add_67879 <= p35_add_67879_comb;
    p35_add_67663 <= p34_add_67663;
    p35_add_67646 <= p34_add_67646;
    p35_add_67487 <= p34_add_67487;
    p35_add_67470 <= p34_add_67470;
    p35_add_67453 <= p34_add_67453;
    p35_add_67780 <= p34_add_67780;
    p35_add_67283 <= p34_add_67283;
    p35_add_67629 <= p34_add_67629;
    p35_add_67249 <= p34_add_67249;
    p35_add_67611 <= p34_add_67611;
    p35_add_67232 <= p34_add_67232;
    p35_add_67436 <= p34_add_67436;
    p35_add_67038 <= p34_add_67038;
    p35_add_67418 <= p34_add_67418;
    p35_add_66118 <= p34_add_66118;
    p35_add_67214 <= p34_add_67214;
  end

  // ===== Pipe stage 36:
  wire [31:0] p36_add_67930_comb;
  wire [31:0] p36_and_67972_comb;
  wire [31:0] p36_add_67952_comb;
  wire [31:0] p36_add_67954_comb;
  wire [31:0] p36_add_67976_comb;
  wire [31:0] p36_add_67955_comb;
  wire [31:0] p36_add_67977_comb;
  assign p36_add_67930_comb = p35_add_67400 + p35_add_67856;
  assign p36_and_67972_comb = p35_add_67879 & p35_add_67762;
  assign p36_add_67952_comb = {p36_add_67930_comb[5:0] ^ p36_add_67930_comb[10:5] ^ p36_add_67930_comb[24:19], p36_add_67930_comb[31:27] ^ p36_add_67930_comb[4:0] ^ p36_add_67930_comb[18:14], p36_add_67930_comb[26:13] ^ p36_add_67930_comb[31:18] ^ p36_add_67930_comb[13:0], p36_add_67930_comb[12:6] ^ p36_add_67930_comb[17:11] ^ p36_add_67930_comb[31:25]} + (p36_add_67930_comb & p35_add_67831 ^ ~(p36_add_67930_comb | ~p35_add_67714));
  assign p36_add_67954_comb = p36_add_67952_comb + 32'ha81a_664b;
  assign p36_add_67976_comb = {p35_add_67879[1:0] ^ p35_add_67879[12:11] ^ p35_add_67879[21:20], p35_add_67879[31:21] ^ p35_add_67879[10:0] ^ p35_add_67879[19:9], p35_add_67879[20:12] ^ p35_add_67879[31:23] ^ p35_add_67879[8:0], p35_add_67879[11:2] ^ p35_add_67879[22:13] ^ p35_add_67879[31:22]} + (p36_and_67972_comb ^ p35_add_67879 & p35_add_67593 ^ p35_and_67874);
  assign p36_add_67955_comb = p36_add_67954_comb + p35_add_67857;
  assign p36_add_67977_comb = p35_add_67856 + p36_add_67976_comb;

  // Registers for pipe stage 36:
  reg [31:0] p36_add_67714;
  reg [31:0] p36_add_67831;
  reg [31:0] p36_add_67930;
  reg [31:0] p36_add_67593;
  reg [31:0] p36_add_67955;
  reg [31:0] p36_add_67762;
  reg [31:0] p36_add_67879;
  reg [31:0] p36_and_67972;
  reg [31:0] p36_add_67977;
  reg [31:0] p36_add_67663;
  reg [31:0] p36_add_67646;
  reg [31:0] p36_add_67487;
  reg [31:0] p36_add_67470;
  reg [31:0] p36_add_67453;
  reg [31:0] p36_add_67780;
  reg [31:0] p36_add_67283;
  reg [31:0] p36_add_67629;
  reg [31:0] p36_add_67249;
  reg [31:0] p36_add_67611;
  reg [31:0] p36_add_67232;
  reg [31:0] p36_add_67436;
  reg [31:0] p36_add_67038;
  reg [31:0] p36_add_67418;
  reg [31:0] p36_add_66118;
  reg [31:0] p36_add_67214;
  always_ff @ (posedge clk) begin
    p36_add_67714 <= p35_add_67714;
    p36_add_67831 <= p35_add_67831;
    p36_add_67930 <= p36_add_67930_comb;
    p36_add_67593 <= p35_add_67593;
    p36_add_67955 <= p36_add_67955_comb;
    p36_add_67762 <= p35_add_67762;
    p36_add_67879 <= p35_add_67879;
    p36_and_67972 <= p36_and_67972_comb;
    p36_add_67977 <= p36_add_67977_comb;
    p36_add_67663 <= p35_add_67663;
    p36_add_67646 <= p35_add_67646;
    p36_add_67487 <= p35_add_67487;
    p36_add_67470 <= p35_add_67470;
    p36_add_67453 <= p35_add_67453;
    p36_add_67780 <= p35_add_67780;
    p36_add_67283 <= p35_add_67283;
    p36_add_67629 <= p35_add_67629;
    p36_add_67249 <= p35_add_67249;
    p36_add_67611 <= p35_add_67611;
    p36_add_67232 <= p35_add_67232;
    p36_add_67436 <= p35_add_67436;
    p36_add_67038 <= p35_add_67038;
    p36_add_67418 <= p35_add_67418;
    p36_add_66118 <= p35_add_66118;
    p36_add_67214 <= p35_add_67214;
  end

  // ===== Pipe stage 37:
  wire [1:0] p37_bit_slice_68078_comb;
  wire [31:0] p37_and_68076_comb;
  wire [31:0] p37_add_68028_comb;
  wire [31:0] p37_add_68081_comb;
  wire [31:0] p37_add_68120_comb;
  wire [31:0] p37_add_68082_comb;
  wire [31:0] p37_add_68121_comb;
  wire [27:0] p37_add_68050_comb;
  wire [31:0] p37_and_68099_comb;
  wire [31:0] p37_add_68055_comb;
  wire [31:0] p37_add_68056_comb;
  wire [31:0] p37_add_68057_comb;
  wire [31:0] p37_add_68117_comb;
  wire [31:0] p37_add_68138_comb;
  wire [31:0] p37_add_68058_comb;
  wire [31:0] p37_add_68059_comb;
  wire [31:0] p37_add_68119_comb;
  wire [31:0] p37_add_68206_comb;
  wire [31:0] p37_add_68189_comb;
  wire [31:0] p37_add_68172_comb;
  wire [31:0] p37_add_68156_comb;
  wire [31:0] p37_add_68139_comb;
  assign p37_bit_slice_68078_comb = p36_add_67232[1:0];
  assign p37_and_68076_comb = p36_add_67977 & p36_add_67879;
  assign p37_add_68028_comb = p36_add_67593 + p36_add_67955;
  assign p37_add_68081_comb = {p36_add_67977[1:0] ^ p36_add_67977[12:11] ^ p36_add_67977[21:20], p36_add_67977[31:21] ^ p36_add_67977[10:0] ^ p36_add_67977[19:9], p36_add_67977[20:12] ^ p36_add_67977[31:23] ^ p36_add_67977[8:0], p36_add_67977[11:2] ^ p36_add_67977[22:13] ^ p36_add_67977[31:22]} + (p37_and_68076_comb ^ p36_add_67977 & p36_add_67762 ^ p36_and_67972);
  assign p37_add_68120_comb = p36_add_67214 + {p36_add_67232[16:7] ^ p36_add_67232[18:9], p36_add_67232[6:0] ^ p36_add_67232[8:2] ^ p36_add_67232[31:25], p36_add_67232[31:30] ^ p37_bit_slice_68078_comb ^ p36_add_67232[24:23], p36_add_67232[29:17] ^ p36_add_67232[31:19] ^ p36_add_67232[22:10]};
  assign p37_add_68082_comb = p36_add_67955 + p37_add_68081_comb;
  assign p37_add_68121_comb = p36_add_67249 + p37_add_68120_comb;
  assign p37_add_68050_comb = p36_add_67418[31:4] + 28'hc24_b8b7;
  assign p37_and_68099_comb = p37_add_68082_comb & p36_add_67977;
  assign p37_add_68055_comb = {p37_add_68028_comb[5:0] ^ p37_add_68028_comb[10:5] ^ p37_add_68028_comb[24:19], p37_add_68028_comb[31:27] ^ p37_add_68028_comb[4:0] ^ p37_add_68028_comb[18:14], p37_add_68028_comb[26:13] ^ p37_add_68028_comb[31:18] ^ p37_add_68028_comb[13:0], p37_add_68028_comb[12:6] ^ p37_add_68028_comb[17:11] ^ p37_add_68028_comb[31:25]} + p36_add_67714;
  assign p37_add_68056_comb = (p37_add_68028_comb & p36_add_67930 ^ ~(p37_add_68028_comb | ~p36_add_67831)) + {p37_add_68050_comb, p36_add_67418[3:0]};
  assign p37_add_68057_comb = p37_add_68055_comb + p37_add_68056_comb;
  assign p37_add_68117_comb = {p37_add_68082_comb[1:0] ^ p37_add_68082_comb[12:11] ^ p37_add_68082_comb[21:20], p37_add_68082_comb[31:21] ^ p37_add_68082_comb[10:0] ^ p37_add_68082_comb[19:9], p37_add_68082_comb[20:12] ^ p37_add_68082_comb[31:23] ^ p37_add_68082_comb[8:0], p37_add_68082_comb[11:2] ^ p37_add_68082_comb[22:13] ^ p37_add_68082_comb[31:22]} + (p37_and_68099_comb ^ p37_add_68082_comb & p36_add_67879 ^ p37_and_68076_comb);
  assign p37_add_68138_comb = p36_add_67418 + {p37_add_68121_comb[16:7] ^ p37_add_68121_comb[18:9], p37_add_68121_comb[6:0] ^ p37_add_68121_comb[8:2] ^ p37_add_68121_comb[31:25], p37_add_68121_comb[31:30] ^ p37_add_68121_comb[1:0] ^ p37_add_68121_comb[24:23], p37_add_68121_comb[29:17] ^ p37_add_68121_comb[31:19] ^ p37_add_68121_comb[22:10]};
  assign p37_add_68058_comb = p36_add_67762 + p37_add_68057_comb;
  assign p37_add_68059_comb = p36_add_67831 + p36_add_67038;
  assign p37_add_68119_comb = p37_add_68057_comb + p37_add_68117_comb;
  assign p37_add_68206_comb = {p36_add_67436[6:4] ^ p36_add_67436[17:15], p36_add_67436[3:0] ^ p36_add_67436[14:11] ^ p36_add_67436[31:28], p36_add_67436[31:21] ^ p36_add_67436[10:0] ^ p36_add_67436[27:17], p36_add_67436[20:7] ^ p36_add_67436[31:18] ^ p36_add_67436[16:3]} + p36_add_67038;
  assign p37_add_68189_comb = {p36_add_67038[6:4] ^ p36_add_67038[17:15], p36_add_67038[3:0] ^ p36_add_67038[14:11] ^ p36_add_67038[31:28], p36_add_67038[31:21] ^ p36_add_67038[10:0] ^ p36_add_67038[27:17], p36_add_67038[20:7] ^ p36_add_67038[31:18] ^ p36_add_67038[16:3]} + p36_add_67418;
  assign p37_add_68172_comb = {p36_add_67418[6:4] ^ p36_add_67418[17:15], p36_add_67418[3:0] ^ p36_add_67418[14:11] ^ p36_add_67418[31:28], p36_add_67418[31:21] ^ p36_add_67418[10:0] ^ p36_add_67418[27:17], p36_add_67418[20:7] ^ p36_add_67418[31:18] ^ p36_add_67418[16:3]} + p36_add_66118;
  assign p37_add_68156_comb = {p36_add_66118[6:4] ^ p36_add_66118[17:15], p36_add_66118[3:0] ^ p36_add_66118[14:11] ^ p36_add_66118[31:28], p36_add_66118[31:21] ^ p36_add_66118[10:0] ^ p36_add_66118[27:17], p36_add_66118[20:7] ^ p36_add_66118[31:18] ^ p36_add_66118[16:3]} + p36_add_67214;
  assign p37_add_68139_comb = p36_add_67283 + p37_add_68138_comb;

  // Registers for pipe stage 37:
  reg [31:0] p37_add_67930;
  reg [31:0] p37_add_68028;
  reg [31:0] p37_add_68058;
  reg [31:0] p37_add_68059;
  reg [31:0] p37_add_67879;
  reg [31:0] p37_add_67977;
  reg [1:0] p37_bit_slice_68078;
  reg [31:0] p37_add_68082;
  reg [31:0] p37_and_68099;
  reg [31:0] p37_add_68119;
  reg [31:0] p37_add_68206;
  reg [31:0] p37_add_68189;
  reg [31:0] p37_add_68172;
  reg [31:0] p37_add_68156;
  reg [31:0] p37_add_67663;
  reg [31:0] p37_add_67646;
  reg [31:0] p37_add_67487;
  reg [31:0] p37_add_67470;
  reg [31:0] p37_add_67453;
  reg [31:0] p37_add_67780;
  reg [31:0] p37_add_68139;
  reg [31:0] p37_add_67629;
  reg [31:0] p37_add_68121;
  reg [31:0] p37_add_67611;
  reg [31:0] p37_add_67232;
  reg [31:0] p37_add_67436;
  always_ff @ (posedge clk) begin
    p37_add_67930 <= p36_add_67930;
    p37_add_68028 <= p37_add_68028_comb;
    p37_add_68058 <= p37_add_68058_comb;
    p37_add_68059 <= p37_add_68059_comb;
    p37_add_67879 <= p36_add_67879;
    p37_add_67977 <= p36_add_67977;
    p37_bit_slice_68078 <= p37_bit_slice_68078_comb;
    p37_add_68082 <= p37_add_68082_comb;
    p37_and_68099 <= p37_and_68099_comb;
    p37_add_68119 <= p37_add_68119_comb;
    p37_add_68206 <= p37_add_68206_comb;
    p37_add_68189 <= p37_add_68189_comb;
    p37_add_68172 <= p37_add_68172_comb;
    p37_add_68156 <= p37_add_68156_comb;
    p37_add_67663 <= p36_add_67663;
    p37_add_67646 <= p36_add_67646;
    p37_add_67487 <= p36_add_67487;
    p37_add_67470 <= p36_add_67470;
    p37_add_67453 <= p36_add_67453;
    p37_add_67780 <= p36_add_67780;
    p37_add_68139 <= p37_add_68139_comb;
    p37_add_67629 <= p36_add_67629;
    p37_add_68121 <= p37_add_68121_comb;
    p37_add_67611 <= p36_add_67611;
    p37_add_67232 <= p36_add_67232;
    p37_add_67436 <= p36_add_67436;
  end

  // ===== Pipe stage 38:
  wire [31:0] p38_add_68324_comb;
  wire [31:0] p38_add_68325_comb;
  wire [31:0] p38_add_68280_comb;
  wire [31:0] p38_and_68302_comb;
  wire [31:0] p38_add_68282_comb;
  wire [31:0] p38_add_68283_comb;
  wire [31:0] p38_add_68306_comb;
  wire [31:0] p38_add_68342_comb;
  wire [31:0] p38_add_68284_comb;
  wire [31:0] p38_add_68285_comb;
  wire [31:0] p38_add_68307_comb;
  wire [31:0] p38_add_68360_comb;
  wire [31:0] p38_add_68343_comb;
  assign p38_add_68324_comb = p37_add_67436 + {p37_add_68139[16:7] ^ p37_add_68139[18:9], p37_add_68139[6:0] ^ p37_add_68139[8:2] ^ p37_add_68139[31:25], p37_add_68139[31:30] ^ p37_add_68139[1:0] ^ p37_add_68139[24:23], p37_add_68139[29:17] ^ p37_add_68139[31:19] ^ p37_add_68139[22:10]};
  assign p38_add_68325_comb = p37_add_67453 + p38_add_68324_comb;
  assign p38_add_68280_comb = {p37_add_68058[5:0] ^ p37_add_68058[10:5] ^ p37_add_68058[24:19], p37_add_68058[31:27] ^ p37_add_68058[4:0] ^ p37_add_68058[18:14], p37_add_68058[26:13] ^ p37_add_68058[31:18] ^ p37_add_68058[13:0], p37_add_68058[12:6] ^ p37_add_68058[17:11] ^ p37_add_68058[31:25]} + (p37_add_68058 & p37_add_68028 ^ ~(p37_add_68058 | ~p37_add_67930));
  assign p38_and_68302_comb = p37_add_68119 & p37_add_68082;
  assign p38_add_68282_comb = p38_add_68280_comb + 32'hc76c_51a3;
  assign p38_add_68283_comb = p38_add_68282_comb + p37_add_68059;
  assign p38_add_68306_comb = {p37_add_68119[1:0] ^ p37_add_68119[12:11] ^ p37_add_68119[21:20], p37_add_68119[31:21] ^ p37_add_68119[10:0] ^ p37_add_68119[19:9], p37_add_68119[20:12] ^ p37_add_68119[31:23] ^ p37_add_68119[8:0], p37_add_68119[11:2] ^ p37_add_68119[22:13] ^ p37_add_68119[31:22]} + (p38_and_68302_comb ^ p37_add_68119 & p37_add_67977 ^ p37_and_68099);
  assign p38_add_68342_comb = p37_add_67611 + {p38_add_68325_comb[16:7] ^ p38_add_68325_comb[18:9], p38_add_68325_comb[6:0] ^ p38_add_68325_comb[8:2] ^ p38_add_68325_comb[31:25], p38_add_68325_comb[31:30] ^ p38_add_68325_comb[1:0] ^ p38_add_68325_comb[24:23], p38_add_68325_comb[29:17] ^ p38_add_68325_comb[31:19] ^ p38_add_68325_comb[22:10]};
  assign p38_add_68284_comb = p37_add_67879 + p38_add_68283_comb;
  assign p38_add_68285_comb = p37_add_67930 + p37_add_67436;
  assign p38_add_68307_comb = p38_add_68283_comb + p38_add_68306_comb;
  assign p38_add_68360_comb = {p37_add_67232[6:4] ^ p37_add_67232[17:15], p37_add_67232[3:0] ^ p37_add_67232[14:11] ^ p37_add_67232[31:28], p37_add_67232[31:21] ^ p37_add_67232[10:0] ^ p37_add_67232[27:17], p37_add_67232[20:7] ^ p37_add_67232[31:18] ^ p37_add_67232[16:3]} + p37_add_67436;
  assign p38_add_68343_comb = p37_add_67487 + p38_add_68342_comb;

  // Registers for pipe stage 38:
  reg [31:0] p38_add_68028;
  reg [31:0] p38_add_68058;
  reg [31:0] p38_add_68284;
  reg [31:0] p38_add_68285;
  reg [31:0] p38_add_67977;
  reg [1:0] p38_bit_slice_68078;
  reg [31:0] p38_add_68082;
  reg [31:0] p38_add_68119;
  reg [31:0] p38_and_68302;
  reg [31:0] p38_add_68307;
  reg [31:0] p38_add_68360;
  reg [31:0] p38_add_68206;
  reg [31:0] p38_add_68189;
  reg [31:0] p38_add_68172;
  reg [31:0] p38_add_68156;
  reg [31:0] p38_add_67663;
  reg [31:0] p38_add_67646;
  reg [31:0] p38_add_68343;
  reg [31:0] p38_add_67470;
  reg [31:0] p38_add_68325;
  reg [31:0] p38_add_67780;
  reg [31:0] p38_add_68139;
  reg [31:0] p38_add_67629;
  reg [31:0] p38_add_68121;
  reg [31:0] p38_add_67611;
  reg [31:0] p38_add_67232;
  always_ff @ (posedge clk) begin
    p38_add_68028 <= p37_add_68028;
    p38_add_68058 <= p37_add_68058;
    p38_add_68284 <= p38_add_68284_comb;
    p38_add_68285 <= p38_add_68285_comb;
    p38_add_67977 <= p37_add_67977;
    p38_bit_slice_68078 <= p37_bit_slice_68078;
    p38_add_68082 <= p37_add_68082;
    p38_add_68119 <= p37_add_68119;
    p38_and_68302 <= p38_and_68302_comb;
    p38_add_68307 <= p38_add_68307_comb;
    p38_add_68360 <= p38_add_68360_comb;
    p38_add_68206 <= p37_add_68206;
    p38_add_68189 <= p37_add_68189;
    p38_add_68172 <= p37_add_68172;
    p38_add_68156 <= p37_add_68156;
    p38_add_67663 <= p37_add_67663;
    p38_add_67646 <= p37_add_67646;
    p38_add_68343 <= p38_add_68343_comb;
    p38_add_67470 <= p37_add_67470;
    p38_add_68325 <= p38_add_68325_comb;
    p38_add_67780 <= p37_add_67780;
    p38_add_68139 <= p37_add_68139;
    p38_add_67629 <= p37_add_67629;
    p38_add_68121 <= p37_add_68121;
    p38_add_67611 <= p37_add_67611;
    p38_add_67232 <= p37_add_67232;
  end

  // ===== Pipe stage 39:
  wire [31:0] p39_add_68521_comb;
  wire [31:0] p39_add_68485_comb;
  wire [31:0] p39_add_68522_comb;
  wire [31:0] p39_add_68486_comb;
  wire [31:0] p39_add_68434_comb;
  wire [31:0] p39_and_68459_comb;
  wire [31:0] p39_add_68436_comb;
  wire [31:0] p39_add_68437_comb;
  wire [29:0] p39_add_68441_comb;
  wire [31:0] p39_add_68463_comb;
  wire [29:0] p39_add_68467_comb;
  wire [31:0] p39_add_68539_comb;
  wire [31:0] p39_add_68503_comb;
  wire [31:0] p39_add_68438_comb;
  wire [31:0] p39_concat_68442_comb;
  wire [31:0] p39_add_68464_comb;
  wire [31:0] p39_concat_68469_comb;
  wire [31:0] p39_add_68557_comb;
  wire [31:0] p39_add_68540_comb;
  wire [31:0] p39_add_68504_comb;
  assign p39_add_68521_comb = p38_add_67629 + {p38_add_68343[16:7] ^ p38_add_68343[18:9], p38_add_68343[6:0] ^ p38_add_68343[8:2] ^ p38_add_68343[31:25], p38_add_68343[31:30] ^ p38_add_68343[1:0] ^ p38_add_68343[24:23], p38_add_68343[29:17] ^ p38_add_68343[31:19] ^ p38_add_68343[22:10]};
  assign p39_add_68485_comb = p38_add_67232 + {p38_add_67780[16:7] ^ p38_add_67780[18:9], p38_add_67780[6:0] ^ p38_add_67780[8:2] ^ p38_add_67780[31:25], p38_add_67780[31:30] ^ p38_add_67780[1:0] ^ p38_add_67780[24:23], p38_add_67780[29:17] ^ p38_add_67780[31:19] ^ p38_add_67780[22:10]};
  assign p39_add_68522_comb = p38_add_67663 + p39_add_68521_comb;
  assign p39_add_68486_comb = p38_add_67470 + p39_add_68485_comb;
  assign p39_add_68434_comb = {p38_add_68284[5:0] ^ p38_add_68284[10:5] ^ p38_add_68284[24:19], p38_add_68284[31:27] ^ p38_add_68284[4:0] ^ p38_add_68284[18:14], p38_add_68284[26:13] ^ p38_add_68284[31:18] ^ p38_add_68284[13:0], p38_add_68284[12:6] ^ p38_add_68284[17:11] ^ p38_add_68284[31:25]} + (p38_add_68284 & p38_add_68058 ^ ~(p38_add_68284 | ~p38_add_68028));
  assign p39_and_68459_comb = p38_add_68307 & p38_add_68119;
  assign p39_add_68436_comb = p39_add_68434_comb + 32'hd192_e819;
  assign p39_add_68437_comb = p39_add_68436_comb + p38_add_68285;
  assign p39_add_68441_comb = p38_add_67232[31:2] + 30'h35a6_4189;
  assign p39_add_68463_comb = {p38_add_68307[1:0] ^ p38_add_68307[12:11] ^ p38_add_68307[21:20], p38_add_68307[31:21] ^ p38_add_68307[10:0] ^ p38_add_68307[19:9], p38_add_68307[20:12] ^ p38_add_68307[31:23] ^ p38_add_68307[8:0], p38_add_68307[11:2] ^ p38_add_68307[22:13] ^ p38_add_68307[31:22]} + (p39_and_68459_comb ^ p38_add_68307 & p38_add_68082 ^ p38_and_68302);
  assign p39_add_68467_comb = p38_add_67780[31:2] + 30'h09d2_1dd3;
  assign p39_add_68539_comb = p38_add_67780 + {p39_add_68522_comb[16:7] ^ p39_add_68522_comb[18:9], p39_add_68522_comb[6:0] ^ p39_add_68522_comb[8:2] ^ p39_add_68522_comb[31:25], p39_add_68522_comb[31:30] ^ p39_add_68522_comb[1:0] ^ p39_add_68522_comb[24:23], p39_add_68522_comb[29:17] ^ p39_add_68522_comb[31:19] ^ p39_add_68522_comb[22:10]};
  assign p39_add_68503_comb = p38_add_68121 + {p39_add_68486_comb[16:7] ^ p39_add_68486_comb[18:9], p39_add_68486_comb[6:0] ^ p39_add_68486_comb[8:2] ^ p39_add_68486_comb[31:25], p39_add_68486_comb[31:30] ^ p39_add_68486_comb[1:0] ^ p39_add_68486_comb[24:23], p39_add_68486_comb[29:17] ^ p39_add_68486_comb[31:19] ^ p39_add_68486_comb[22:10]};
  assign p39_add_68438_comb = p38_add_67977 + p39_add_68437_comb;
  assign p39_concat_68442_comb = {p39_add_68441_comb, p38_bit_slice_68078};
  assign p39_add_68464_comb = p39_add_68437_comb + p39_add_68463_comb;
  assign p39_concat_68469_comb = {p39_add_68467_comb, p38_add_67780[1:0]};
  assign p39_add_68557_comb = {p38_add_67611[6:4] ^ p38_add_67611[17:15], p38_add_67611[3:0] ^ p38_add_67611[14:11] ^ p38_add_67611[31:28], p38_add_67611[31:21] ^ p38_add_67611[10:0] ^ p38_add_67611[27:17], p38_add_67611[20:7] ^ p38_add_67611[31:18] ^ p38_add_67611[16:3]} + p38_add_67232;
  assign p39_add_68540_comb = p38_add_68172 + p39_add_68539_comb;
  assign p39_add_68504_comb = p38_add_67646 + p39_add_68503_comb;

  // Registers for pipe stage 39:
  reg [31:0] p39_add_68028;
  reg [31:0] p39_add_68058;
  reg [31:0] p39_add_68284;
  reg [31:0] p39_add_68438;
  reg [31:0] p39_concat_68442;
  reg [31:0] p39_add_68082;
  reg [31:0] p39_add_68119;
  reg [31:0] p39_add_68307;
  reg [31:0] p39_and_68459;
  reg [31:0] p39_add_68464;
  reg [31:0] p39_concat_68469;
  reg [31:0] p39_add_68557;
  reg [31:0] p39_add_68360;
  reg [31:0] p39_add_68206;
  reg [31:0] p39_add_68189;
  reg [31:0] p39_add_68540;
  reg [31:0] p39_add_68156;
  reg [31:0] p39_add_68522;
  reg [31:0] p39_add_68504;
  reg [31:0] p39_add_68343;
  reg [31:0] p39_add_68486;
  reg [31:0] p39_add_68325;
  reg [31:0] p39_add_68139;
  reg [31:0] p39_add_67629;
  reg [31:0] p39_add_68121;
  reg [31:0] p39_add_67611;
  always_ff @ (posedge clk) begin
    p39_add_68028 <= p38_add_68028;
    p39_add_68058 <= p38_add_68058;
    p39_add_68284 <= p38_add_68284;
    p39_add_68438 <= p39_add_68438_comb;
    p39_concat_68442 <= p39_concat_68442_comb;
    p39_add_68082 <= p38_add_68082;
    p39_add_68119 <= p38_add_68119;
    p39_add_68307 <= p38_add_68307;
    p39_and_68459 <= p39_and_68459_comb;
    p39_add_68464 <= p39_add_68464_comb;
    p39_concat_68469 <= p39_concat_68469_comb;
    p39_add_68557 <= p39_add_68557_comb;
    p39_add_68360 <= p38_add_68360;
    p39_add_68206 <= p38_add_68206;
    p39_add_68189 <= p38_add_68189;
    p39_add_68540 <= p39_add_68540_comb;
    p39_add_68156 <= p38_add_68156;
    p39_add_68522 <= p39_add_68522_comb;
    p39_add_68504 <= p39_add_68504_comb;
    p39_add_68343 <= p38_add_68343;
    p39_add_68486 <= p39_add_68486_comb;
    p39_add_68325 <= p38_add_68325;
    p39_add_68139 <= p38_add_68139;
    p39_add_67629 <= p38_add_67629;
    p39_add_68121 <= p38_add_68121;
    p39_add_67611 <= p38_add_67611;
  end

  // ===== Pipe stage 40:
  wire [31:0] p40_add_68631_comb;
  wire [31:0] p40_add_68632_comb;
  wire [31:0] p40_add_68737_comb;
  wire [31:0] p40_add_68701_comb;
  wire [31:0] p40_add_68633_comb;
  wire [31:0] p40_add_68738_comb;
  wire [31:0] p40_add_68702_comb;
  wire [31:0] p40_add_68634_comb;
  wire [31:0] p40_and_68676_comb;
  wire [28:0] p40_add_68678_comb;
  wire [31:0] p40_add_68683_comb;
  wire [28:0] p40_add_68741_comb;
  wire [31:0] p40_add_68760_comb;
  wire [31:0] p40_add_68719_comb;
  wire [31:0] p40_add_68656_comb;
  wire [31:0] p40_add_68657_comb;
  wire [31:0] p40_concat_68682_comb;
  wire [31:0] p40_add_68684_comb;
  wire [31:0] p40_concat_68743_comb;
  wire [31:0] p40_add_68761_comb;
  wire [31:0] p40_add_68720_comb;
  assign p40_add_68631_comb = {p39_add_68438[5:0] ^ p39_add_68438[10:5] ^ p39_add_68438[24:19], p39_add_68438[31:27] ^ p39_add_68438[4:0] ^ p39_add_68438[18:14], p39_add_68438[26:13] ^ p39_add_68438[31:18] ^ p39_add_68438[13:0], p39_add_68438[12:6] ^ p39_add_68438[17:11] ^ p39_add_68438[31:25]} + p39_add_68028;
  assign p40_add_68632_comb = (p39_add_68438 & p39_add_68284 ^ ~(p39_add_68438 | ~p39_add_68058)) + p39_concat_68442;
  assign p40_add_68737_comb = p39_add_68486 + {p39_add_68540[16:7] ^ p39_add_68540[18:9], p39_add_68540[6:0] ^ p39_add_68540[8:2] ^ p39_add_68540[31:25], p39_add_68540[31:30] ^ p39_add_68540[1:0] ^ p39_add_68540[24:23], p39_add_68540[29:17] ^ p39_add_68540[31:19] ^ p39_add_68540[22:10]};
  assign p40_add_68701_comb = p39_add_68139 + {p39_add_68504[16:7] ^ p39_add_68504[18:9], p39_add_68504[6:0] ^ p39_add_68504[8:2] ^ p39_add_68504[31:25], p39_add_68504[31:30] ^ p39_add_68504[1:0] ^ p39_add_68504[24:23], p39_add_68504[29:17] ^ p39_add_68504[31:19] ^ p39_add_68504[22:10]};
  assign p40_add_68633_comb = p40_add_68631_comb + p40_add_68632_comb;
  assign p40_add_68738_comb = p39_add_68206 + p40_add_68737_comb;
  assign p40_add_68702_comb = p39_add_68156 + p40_add_68701_comb;
  assign p40_add_68634_comb = p39_add_68082 + p40_add_68633_comb;
  assign p40_and_68676_comb = p39_add_68464 & p39_add_68307;
  assign p40_add_68678_comb = p39_add_68139[31:3] + 29'h03c6_ed81;
  assign p40_add_68683_comb = {p39_add_68464[1:0] ^ p39_add_68464[12:11] ^ p39_add_68464[21:20], p39_add_68464[31:21] ^ p39_add_68464[10:0] ^ p39_add_68464[19:9], p39_add_68464[20:12] ^ p39_add_68464[31:23] ^ p39_add_68464[8:0], p39_add_68464[11:2] ^ p39_add_68464[22:13] ^ p39_add_68464[31:22]} + (p40_and_68676_comb ^ p39_add_68464 & p39_add_68119 ^ p39_and_68459);
  assign p40_add_68741_comb = p40_add_68738_comb[31:3] + 29'h1198_e041;
  assign p40_add_68760_comb = p39_add_68504 + {p40_add_68738_comb[16:7] ^ p40_add_68738_comb[18:9], p40_add_68738_comb[6:0] ^ p40_add_68738_comb[8:2] ^ p40_add_68738_comb[31:25], p40_add_68738_comb[31:30] ^ p40_add_68738_comb[1:0] ^ p40_add_68738_comb[24:23], p40_add_68738_comb[29:17] ^ p40_add_68738_comb[31:19] ^ p40_add_68738_comb[22:10]};
  assign p40_add_68719_comb = p39_add_68325 + {p40_add_68702_comb[16:7] ^ p40_add_68702_comb[18:9], p40_add_68702_comb[6:0] ^ p40_add_68702_comb[8:2] ^ p40_add_68702_comb[31:25], p40_add_68702_comb[31:30] ^ p40_add_68702_comb[1:0] ^ p40_add_68702_comb[24:23], p40_add_68702_comb[29:17] ^ p40_add_68702_comb[31:19] ^ p40_add_68702_comb[22:10]};
  assign p40_add_68656_comb = {p40_add_68634_comb[5:0] ^ p40_add_68634_comb[10:5] ^ p40_add_68634_comb[24:19], p40_add_68634_comb[31:27] ^ p40_add_68634_comb[4:0] ^ p40_add_68634_comb[18:14], p40_add_68634_comb[26:13] ^ p40_add_68634_comb[31:18] ^ p40_add_68634_comb[13:0], p40_add_68634_comb[12:6] ^ p40_add_68634_comb[17:11] ^ p40_add_68634_comb[31:25]} + (p40_add_68634_comb & p39_add_68438 ^ ~(p40_add_68634_comb | ~p39_add_68284));
  assign p40_add_68657_comb = p39_add_68058 + p39_add_67611;
  assign p40_concat_68682_comb = {p40_add_68678_comb, p39_add_68139[2:0]};
  assign p40_add_68684_comb = p40_add_68633_comb + p40_add_68683_comb;
  assign p40_concat_68743_comb = {p40_add_68741_comb, p40_add_68738_comb[2:0]};
  assign p40_add_68761_comb = p39_add_68557 + p40_add_68760_comb;
  assign p40_add_68720_comb = p39_add_68189 + p40_add_68719_comb;

  // Registers for pipe stage 40:
  reg [31:0] p40_add_68284;
  reg [31:0] p40_add_68438;
  reg [31:0] p40_add_68634;
  reg [31:0] p40_add_68656;
  reg [31:0] p40_add_68657;
  reg [31:0] p40_add_68119;
  reg [31:0] p40_add_68307;
  reg [31:0] p40_add_68464;
  reg [31:0] p40_and_68676;
  reg [31:0] p40_concat_68682;
  reg [31:0] p40_add_68684;
  reg [31:0] p40_concat_68469;
  reg [31:0] p40_concat_68743;
  reg [31:0] p40_add_68761;
  reg [31:0] p40_add_68360;
  reg [31:0] p40_add_68720;
  reg [31:0] p40_add_68540;
  reg [31:0] p40_add_68702;
  reg [31:0] p40_add_68522;
  reg [31:0] p40_add_68504;
  reg [31:0] p40_add_68343;
  reg [31:0] p40_add_68486;
  reg [31:0] p40_add_68325;
  reg [31:0] p40_add_67629;
  reg [31:0] p40_add_68121;
  reg [31:0] p40_add_67611;
  always_ff @ (posedge clk) begin
    p40_add_68284 <= p39_add_68284;
    p40_add_68438 <= p39_add_68438;
    p40_add_68634 <= p40_add_68634_comb;
    p40_add_68656 <= p40_add_68656_comb;
    p40_add_68657 <= p40_add_68657_comb;
    p40_add_68119 <= p39_add_68119;
    p40_add_68307 <= p39_add_68307;
    p40_add_68464 <= p39_add_68464;
    p40_and_68676 <= p40_and_68676_comb;
    p40_concat_68682 <= p40_concat_68682_comb;
    p40_add_68684 <= p40_add_68684_comb;
    p40_concat_68469 <= p39_concat_68469;
    p40_concat_68743 <= p40_concat_68743_comb;
    p40_add_68761 <= p40_add_68761_comb;
    p40_add_68360 <= p39_add_68360;
    p40_add_68720 <= p40_add_68720_comb;
    p40_add_68540 <= p39_add_68540;
    p40_add_68702 <= p40_add_68702_comb;
    p40_add_68522 <= p39_add_68522;
    p40_add_68504 <= p39_add_68504;
    p40_add_68343 <= p39_add_68343;
    p40_add_68486 <= p39_add_68486;
    p40_add_68325 <= p39_add_68325;
    p40_add_67629 <= p39_add_67629;
    p40_add_68121 <= p39_add_68121;
    p40_add_67611 <= p39_add_67611;
  end

  // ===== Pipe stage 41:
  wire [31:0] p41_add_68815_comb;
  wire [31:0] p41_add_68816_comb;
  wire [31:0] p41_add_68817_comb;
  wire [31:0] p41_and_68862_comb;
  wire [27:0] p41_add_68839_comb;
  wire [31:0] p41_add_68866_comb;
  wire [30:0] p41_add_68870_comb;
  wire [29:0] p41_add_68875_comb;
  wire [31:0] p41_add_68893_comb;
  wire [31:0] p41_add_68867_comb;
  wire [31:0] p41_concat_68872_comb;
  wire [31:0] p41_concat_68877_comb;
  wire [3:0] p41_xor_68897_comb;
  wire [31:0] p41_add_68894_comb;
  wire [31:0] p41_add_68844_comb;
  wire [31:0] p41_add_68845_comb;
  assign p41_add_68815_comb = p40_add_68656 + 32'hf40e_3585;
  assign p41_add_68816_comb = p41_add_68815_comb + p40_add_68657;
  assign p41_add_68817_comb = p40_add_68119 + p41_add_68816_comb;
  assign p41_and_68862_comb = p40_add_68684 & p40_add_68464;
  assign p41_add_68839_comb = p40_add_68121[31:4] + 28'h106_aa07;
  assign p41_add_68866_comb = {p40_add_68684[1:0] ^ p40_add_68684[12:11] ^ p40_add_68684[21:20], p40_add_68684[31:21] ^ p40_add_68684[10:0] ^ p40_add_68684[19:9], p40_add_68684[20:12] ^ p40_add_68684[31:23] ^ p40_add_68684[8:0], p40_add_68684[11:2] ^ p40_add_68684[22:13] ^ p40_add_68684[31:22]} + (p41_and_68862_comb ^ p40_add_68684 & p40_add_68307 ^ p40_and_68676);
  assign p41_add_68870_comb = p40_add_68343[31:1] + 31'h276c_5525;
  assign p41_add_68875_comb = p40_add_68720[31:2] + 30'h2132_1e05;
  assign p41_add_68893_comb = p40_add_68343 + {p40_add_68720[16:7] ^ p40_add_68720[18:9], p40_add_68720[6:0] ^ p40_add_68720[8:2] ^ p40_add_68720[31:25], p40_add_68720[31:30] ^ p40_add_68720[1:0] ^ p40_add_68720[24:23], p40_add_68720[29:17] ^ p40_add_68720[31:19] ^ p40_add_68720[22:10]};
  assign p41_add_68867_comb = p41_add_68816_comb + p41_add_68866_comb;
  assign p41_concat_68872_comb = {p41_add_68870_comb, p40_add_68343[0]};
  assign p41_concat_68877_comb = {p41_add_68875_comb, p40_add_68720[1:0]};
  assign p41_xor_68897_comb = p40_add_68121[3:0] ^ p40_add_68121[14:11] ^ p40_add_68121[31:28];
  assign p41_add_68894_comb = p40_add_68360 + p41_add_68893_comb;
  assign p41_add_68844_comb = {p41_add_68817_comb[5:0] ^ p41_add_68817_comb[10:5] ^ p41_add_68817_comb[24:19], p41_add_68817_comb[31:27] ^ p41_add_68817_comb[4:0] ^ p41_add_68817_comb[18:14], p41_add_68817_comb[26:13] ^ p41_add_68817_comb[31:18] ^ p41_add_68817_comb[13:0], p41_add_68817_comb[12:6] ^ p41_add_68817_comb[17:11] ^ p41_add_68817_comb[31:25]} + p40_add_68284;
  assign p41_add_68845_comb = (p41_add_68817_comb & p40_add_68634 ^ ~(p41_add_68817_comb | ~p40_add_68438)) + {p41_add_68839_comb, p40_add_68121[3:0]};

  // Registers for pipe stage 41:
  reg [31:0] p41_add_68438;
  reg [31:0] p41_add_68634;
  reg [31:0] p41_add_68817;
  reg [31:0] p41_add_68307;
  reg [31:0] p41_add_68464;
  reg [31:0] p41_concat_68682;
  reg [31:0] p41_add_68684;
  reg [31:0] p41_and_68862;
  reg [31:0] p41_concat_68469;
  reg [31:0] p41_add_68867;
  reg [31:0] p41_concat_68872;
  reg [31:0] p41_concat_68877;
  reg [31:0] p41_concat_68743;
  reg [3:0] p41_xor_68897;
  reg [31:0] p41_add_68761;
  reg [31:0] p41_add_68894;
  reg [31:0] p41_add_68540;
  reg [31:0] p41_add_68702;
  reg [31:0] p41_add_68522;
  reg [31:0] p41_add_68504;
  reg [31:0] p41_add_68486;
  reg [31:0] p41_add_68325;
  reg [31:0] p41_add_67629;
  reg [31:0] p41_add_68844;
  reg [31:0] p41_add_68845;
  reg [31:0] p41_add_68121;
  reg [31:0] p41_add_67611;
  always_ff @ (posedge clk) begin
    p41_add_68438 <= p40_add_68438;
    p41_add_68634 <= p40_add_68634;
    p41_add_68817 <= p41_add_68817_comb;
    p41_add_68307 <= p40_add_68307;
    p41_add_68464 <= p40_add_68464;
    p41_concat_68682 <= p40_concat_68682;
    p41_add_68684 <= p40_add_68684;
    p41_and_68862 <= p41_and_68862_comb;
    p41_concat_68469 <= p40_concat_68469;
    p41_add_68867 <= p41_add_68867_comb;
    p41_concat_68872 <= p41_concat_68872_comb;
    p41_concat_68877 <= p41_concat_68877_comb;
    p41_concat_68743 <= p40_concat_68743;
    p41_xor_68897 <= p41_xor_68897_comb;
    p41_add_68761 <= p40_add_68761;
    p41_add_68894 <= p41_add_68894_comb;
    p41_add_68540 <= p40_add_68540;
    p41_add_68702 <= p40_add_68702;
    p41_add_68522 <= p40_add_68522;
    p41_add_68504 <= p40_add_68504;
    p41_add_68486 <= p40_add_68486;
    p41_add_68325 <= p40_add_68325;
    p41_add_67629 <= p40_add_67629;
    p41_add_68844 <= p41_add_68844_comb;
    p41_add_68845 <= p41_add_68845_comb;
    p41_add_68121 <= p40_add_68121;
    p41_add_67611 <= p40_add_67611;
  end

  // ===== Pipe stage 42:
  wire [31:0] p42_add_68952_comb;
  wire [31:0] p42_add_68953_comb;
  wire [31:0] p42_and_68999_comb;
  wire [30:0] p42_add_68975_comb;
  wire [31:0] p42_add_69003_comb;
  wire [31:0] p42_add_68980_comb;
  wire [31:0] p42_add_68981_comb;
  wire [31:0] p42_add_69004_comb;
  wire [31:0] p42_add_69005_comb;
  wire [31:0] p42_concat_69021_comb;
  wire [31:0] p42_add_68982_comb;
  assign p42_add_68952_comb = p41_add_68844 + p41_add_68845;
  assign p42_add_68953_comb = p41_add_68307 + p42_add_68952_comb;
  assign p42_and_68999_comb = p41_add_68867 & p41_add_68684;
  assign p42_add_68975_comb = p41_add_67629[31:1] + 31'h0cd2_608b;
  assign p42_add_69003_comb = {p41_add_68867[1:0] ^ p41_add_68867[12:11] ^ p41_add_68867[21:20], p41_add_68867[31:21] ^ p41_add_68867[10:0] ^ p41_add_68867[19:9], p41_add_68867[20:12] ^ p41_add_68867[31:23] ^ p41_add_68867[8:0], p41_add_68867[11:2] ^ p41_add_68867[22:13] ^ p41_add_68867[31:22]} + (p42_and_68999_comb ^ p41_add_68867 & p41_add_68464 ^ p41_and_68862);
  assign p42_add_68980_comb = {p42_add_68953_comb[5:0] ^ p42_add_68953_comb[10:5] ^ p42_add_68953_comb[24:19], p42_add_68953_comb[31:27] ^ p42_add_68953_comb[4:0] ^ p42_add_68953_comb[18:14], p42_add_68953_comb[26:13] ^ p42_add_68953_comb[31:18] ^ p42_add_68953_comb[13:0], p42_add_68953_comb[12:6] ^ p42_add_68953_comb[17:11] ^ p42_add_68953_comb[31:25]} + p41_add_68438;
  assign p42_add_68981_comb = (p42_add_68953_comb & p41_add_68817 ^ ~(p42_add_68953_comb | ~p41_add_68634)) + {p42_add_68975_comb, p41_add_67629[0]};
  assign p42_add_69004_comb = p42_add_68953_comb + p41_add_68325;
  assign p42_add_69005_comb = p42_add_68952_comb + p42_add_69003_comb;
  assign p42_concat_69021_comb = {p41_add_67629[6:4] ^ p41_add_67629[17:15], p41_add_67629[3:0] ^ p41_add_67629[14:11] ^ p41_add_67629[31:28], p41_add_67629[31:21] ^ p41_add_67629[10:0] ^ p41_add_67629[27:17], p41_add_67629[20:7] ^ p41_add_67629[31:18] ^ p41_add_67629[16:3]};
  assign p42_add_68982_comb = p42_add_68980_comb + p42_add_68981_comb;

  // Registers for pipe stage 42:
  reg [31:0] p42_add_68634;
  reg [31:0] p42_add_68817;
  reg [31:0] p42_add_68953;
  reg [31:0] p42_add_68464;
  reg [31:0] p42_concat_68682;
  reg [31:0] p42_add_68684;
  reg [31:0] p42_concat_68469;
  reg [31:0] p42_add_68867;
  reg [31:0] p42_and_68999;
  reg [31:0] p42_add_69004;
  reg [31:0] p42_add_69005;
  reg [31:0] p42_concat_68872;
  reg [31:0] p42_concat_68877;
  reg [31:0] p42_concat_68743;
  reg [3:0] p42_xor_68897;
  reg [31:0] p42_concat_69021;
  reg [31:0] p42_add_68761;
  reg [31:0] p42_add_68894;
  reg [31:0] p42_add_68540;
  reg [31:0] p42_add_68702;
  reg [31:0] p42_add_68522;
  reg [31:0] p42_add_68504;
  reg [31:0] p42_add_68486;
  reg [31:0] p42_add_68982;
  reg [31:0] p42_add_68121;
  reg [31:0] p42_add_67611;
  always_ff @ (posedge clk) begin
    p42_add_68634 <= p41_add_68634;
    p42_add_68817 <= p41_add_68817;
    p42_add_68953 <= p42_add_68953_comb;
    p42_add_68464 <= p41_add_68464;
    p42_concat_68682 <= p41_concat_68682;
    p42_add_68684 <= p41_add_68684;
    p42_concat_68469 <= p41_concat_68469;
    p42_add_68867 <= p41_add_68867;
    p42_and_68999 <= p42_and_68999_comb;
    p42_add_69004 <= p42_add_69004_comb;
    p42_add_69005 <= p42_add_69005_comb;
    p42_concat_68872 <= p41_concat_68872;
    p42_concat_68877 <= p41_concat_68877;
    p42_concat_68743 <= p41_concat_68743;
    p42_xor_68897 <= p41_xor_68897;
    p42_concat_69021 <= p42_concat_69021_comb;
    p42_add_68761 <= p41_add_68761;
    p42_add_68894 <= p41_add_68894;
    p42_add_68540 <= p41_add_68540;
    p42_add_68702 <= p41_add_68702;
    p42_add_68522 <= p41_add_68522;
    p42_add_68504 <= p41_add_68504;
    p42_add_68486 <= p41_add_68486;
    p42_add_68982 <= p42_add_68982_comb;
    p42_add_68121 <= p41_add_68121;
    p42_add_67611 <= p41_add_67611;
  end

  // ===== Pipe stage 43:
  wire [31:0] p43_add_69074_comb;
  wire [31:0] p43_and_69121_comb;
  wire [31:0] p43_add_69125_comb;
  wire [31:0] p43_add_69126_comb;
  wire [31:0] p43_add_69096_comb;
  wire [31:0] p43_add_69097_comb;
  wire [31:0] p43_add_69098_comb;
  wire [31:0] p43_and_69144_comb;
  wire [31:0] p43_add_69099_comb;
  wire [31:0] p43_add_69148_comb;
  wire [31:0] p43_xor_69103_comb;
  wire [31:0] p43_not_69104_comb;
  wire [31:0] p43_add_69127_comb;
  wire [31:0] p43_add_69149_comb;
  assign p43_add_69074_comb = p42_add_68464 + p42_add_68982;
  assign p43_and_69121_comb = p42_add_69005 & p42_add_68867;
  assign p43_add_69125_comb = {p42_add_69005[1:0] ^ p42_add_69005[12:11] ^ p42_add_69005[21:20], p42_add_69005[31:21] ^ p42_add_69005[10:0] ^ p42_add_69005[19:9], p42_add_69005[20:12] ^ p42_add_69005[31:23] ^ p42_add_69005[8:0], p42_add_69005[11:2] ^ p42_add_69005[22:13] ^ p42_add_69005[31:22]} + (p43_and_69121_comb ^ p42_add_69005 & p42_add_68684 ^ p42_and_68999);
  assign p43_add_69126_comb = p42_add_68982 + p43_add_69125_comb;
  assign p43_add_69096_comb = {p43_add_69074_comb[5:0] ^ p43_add_69074_comb[10:5] ^ p43_add_69074_comb[24:19], p43_add_69074_comb[31:27] ^ p43_add_69074_comb[4:0] ^ p43_add_69074_comb[18:14], p43_add_69074_comb[26:13] ^ p43_add_69074_comb[31:18] ^ p43_add_69074_comb[13:0], p43_add_69074_comb[12:6] ^ p43_add_69074_comb[17:11] ^ p43_add_69074_comb[31:25]} + p42_add_68634;
  assign p43_add_69097_comb = (p43_add_69074_comb & p42_add_68953 ^ ~(p43_add_69074_comb | ~p42_add_68817)) + p42_concat_68682;
  assign p43_add_69098_comb = p43_add_69096_comb + p43_add_69097_comb;
  assign p43_and_69144_comb = p43_add_69126_comb & p42_add_69005;
  assign p43_add_69099_comb = p42_add_68684 + p43_add_69098_comb;
  assign p43_add_69148_comb = {p43_add_69126_comb[1:0] ^ p43_add_69126_comb[12:11] ^ p43_add_69126_comb[21:20], p43_add_69126_comb[31:21] ^ p43_add_69126_comb[10:0] ^ p43_add_69126_comb[19:9], p43_add_69126_comb[20:12] ^ p43_add_69126_comb[31:23] ^ p43_add_69126_comb[8:0], p43_add_69126_comb[11:2] ^ p43_add_69126_comb[22:13] ^ p43_add_69126_comb[31:22]} + (p43_and_69144_comb ^ p43_add_69126_comb & p42_add_68867 ^ p43_and_69121_comb);
  assign p43_xor_69103_comb = p43_add_69099_comb & p43_add_69074_comb ^ ~(p43_add_69099_comb | ~p42_add_68953);
  assign p43_not_69104_comb = ~p43_add_69074_comb;
  assign p43_add_69127_comb = p43_add_69074_comb + p42_add_68486;
  assign p43_add_69149_comb = p43_add_69098_comb + p43_add_69148_comb;

  // Registers for pipe stage 43:
  reg [31:0] p43_add_68817;
  reg [31:0] p43_add_69099;
  reg [31:0] p43_xor_69103;
  reg [31:0] p43_concat_68469;
  reg [31:0] p43_add_68867;
  reg [31:0] p43_not_69104;
  reg [31:0] p43_add_69004;
  reg [31:0] p43_add_69005;
  reg [31:0] p43_add_69127;
  reg [31:0] p43_add_69126;
  reg [31:0] p43_and_69144;
  reg [31:0] p43_concat_68872;
  reg [31:0] p43_add_69149;
  reg [31:0] p43_concat_68877;
  reg [31:0] p43_concat_68743;
  reg [3:0] p43_xor_68897;
  reg [31:0] p43_concat_69021;
  reg [31:0] p43_add_68761;
  reg [31:0] p43_add_68894;
  reg [31:0] p43_add_68540;
  reg [31:0] p43_add_68702;
  reg [31:0] p43_add_68522;
  reg [31:0] p43_add_68504;
  reg [31:0] p43_add_68121;
  reg [31:0] p43_add_67611;
  always_ff @ (posedge clk) begin
    p43_add_68817 <= p42_add_68817;
    p43_add_69099 <= p43_add_69099_comb;
    p43_xor_69103 <= p43_xor_69103_comb;
    p43_concat_68469 <= p42_concat_68469;
    p43_add_68867 <= p42_add_68867;
    p43_not_69104 <= p43_not_69104_comb;
    p43_add_69004 <= p42_add_69004;
    p43_add_69005 <= p42_add_69005;
    p43_add_69127 <= p43_add_69127_comb;
    p43_add_69126 <= p43_add_69126_comb;
    p43_and_69144 <= p43_and_69144_comb;
    p43_concat_68872 <= p42_concat_68872;
    p43_add_69149 <= p43_add_69149_comb;
    p43_concat_68877 <= p42_concat_68877;
    p43_concat_68743 <= p42_concat_68743;
    p43_xor_68897 <= p42_xor_68897;
    p43_concat_69021 <= p42_concat_69021;
    p43_add_68761 <= p42_add_68761;
    p43_add_68894 <= p42_add_68894;
    p43_add_68540 <= p42_add_68540;
    p43_add_68702 <= p42_add_68702;
    p43_add_68522 <= p42_add_68522;
    p43_add_68504 <= p42_add_68504;
    p43_add_68121 <= p42_add_68121;
    p43_add_67611 <= p42_add_67611;
  end

  // ===== Pipe stage 44:
  wire [31:0] p44_add_69217_comb;
  wire [31:0] p44_add_69218_comb;
  wire [31:0] p44_add_69219_comb;
  wire [31:0] p44_add_69220_comb;
  wire [31:0] p44_and_69258_comb;
  wire [31:0] p44_add_69262_comb;
  wire [31:0] p44_add_69241_comb;
  wire [31:0] p44_add_69263_comb;
  wire [31:0] p44_add_69264_comb;
  assign p44_add_69217_comb = {p43_add_69099[5:0] ^ p43_add_69099[10:5] ^ p43_add_69099[24:19], p43_add_69099[31:27] ^ p43_add_69099[4:0] ^ p43_add_69099[18:14], p43_add_69099[26:13] ^ p43_add_69099[31:18] ^ p43_add_69099[13:0], p43_add_69099[12:6] ^ p43_add_69099[17:11] ^ p43_add_69099[31:25]} + p43_add_68817;
  assign p44_add_69218_comb = p43_xor_69103 + p43_concat_68469;
  assign p44_add_69219_comb = p44_add_69217_comb + p44_add_69218_comb;
  assign p44_add_69220_comb = p43_add_68867 + p44_add_69219_comb;
  assign p44_and_69258_comb = p43_add_69149 & p43_add_69126;
  assign p44_add_69262_comb = {p43_add_69149[1:0] ^ p43_add_69149[12:11] ^ p43_add_69149[21:20], p43_add_69149[31:21] ^ p43_add_69149[10:0] ^ p43_add_69149[19:9], p43_add_69149[20:12] ^ p43_add_69149[31:23] ^ p43_add_69149[8:0], p43_add_69149[11:2] ^ p43_add_69149[22:13] ^ p43_add_69149[31:22]} + (p44_and_69258_comb ^ p43_add_69149 & p43_add_69005 ^ p43_and_69144);
  assign p44_add_69241_comb = {p44_add_69220_comb[5:0] ^ p44_add_69220_comb[10:5] ^ p44_add_69220_comb[24:19], p44_add_69220_comb[31:27] ^ p44_add_69220_comb[4:0] ^ p44_add_69220_comb[18:14], p44_add_69220_comb[26:13] ^ p44_add_69220_comb[31:18] ^ p44_add_69220_comb[13:0], p44_add_69220_comb[12:6] ^ p44_add_69220_comb[17:11] ^ p44_add_69220_comb[31:25]} + (p44_add_69220_comb & p43_add_69099 ^ ~(p44_add_69220_comb | p43_not_69104));
  assign p44_add_69263_comb = p44_add_69219_comb + p44_add_69262_comb;
  assign p44_add_69264_comb = p44_add_69220_comb + p43_add_68504;

  // Registers for pipe stage 44:
  reg [31:0] p44_add_69099;
  reg [31:0] p44_add_69220;
  reg [31:0] p44_add_69241;
  reg [31:0] p44_add_69004;
  reg [31:0] p44_add_69005;
  reg [31:0] p44_add_69127;
  reg [31:0] p44_add_69126;
  reg [31:0] p44_concat_68872;
  reg [31:0] p44_add_69149;
  reg [31:0] p44_and_69258;
  reg [31:0] p44_add_69263;
  reg [31:0] p44_add_69264;
  reg [31:0] p44_concat_68877;
  reg [31:0] p44_concat_68743;
  reg [3:0] p44_xor_68897;
  reg [31:0] p44_concat_69021;
  reg [31:0] p44_add_68761;
  reg [31:0] p44_add_68894;
  reg [31:0] p44_add_68540;
  reg [31:0] p44_add_68702;
  reg [31:0] p44_add_68522;
  reg [31:0] p44_add_68121;
  reg [31:0] p44_add_67611;
  always_ff @ (posedge clk) begin
    p44_add_69099 <= p43_add_69099;
    p44_add_69220 <= p44_add_69220_comb;
    p44_add_69241 <= p44_add_69241_comb;
    p44_add_69004 <= p43_add_69004;
    p44_add_69005 <= p43_add_69005;
    p44_add_69127 <= p43_add_69127;
    p44_add_69126 <= p43_add_69126;
    p44_concat_68872 <= p43_concat_68872;
    p44_add_69149 <= p43_add_69149;
    p44_and_69258 <= p44_and_69258_comb;
    p44_add_69263 <= p44_add_69263_comb;
    p44_add_69264 <= p44_add_69264_comb;
    p44_concat_68877 <= p43_concat_68877;
    p44_concat_68743 <= p43_concat_68743;
    p44_xor_68897 <= p43_xor_68897;
    p44_concat_69021 <= p43_concat_69021;
    p44_add_68761 <= p43_add_68761;
    p44_add_68894 <= p43_add_68894;
    p44_add_68540 <= p43_add_68540;
    p44_add_68702 <= p43_add_68702;
    p44_add_68522 <= p43_add_68522;
    p44_add_68121 <= p43_add_68121;
    p44_add_67611 <= p43_add_67611;
  end

  // ===== Pipe stage 45:
  wire [31:0] p45_add_69312_comb;
  wire [31:0] p45_add_69313_comb;
  wire [31:0] p45_add_69314_comb;
  wire [31:0] p45_and_69354_comb;
  wire [31:0] p45_add_69358_comb;
  wire [31:0] p45_add_69336_comb;
  wire [31:0] p45_not_69337_comb;
  wire [31:0] p45_add_69359_comb;
  assign p45_add_69312_comb = p44_add_69241 + 32'h34b0_bcb5;
  assign p45_add_69313_comb = p45_add_69312_comb + p44_add_69004;
  assign p45_add_69314_comb = p44_add_69005 + p45_add_69313_comb;
  assign p45_and_69354_comb = p44_add_69263 & p44_add_69149;
  assign p45_add_69358_comb = {p44_add_69263[1:0] ^ p44_add_69263[12:11] ^ p44_add_69263[21:20], p44_add_69263[31:21] ^ p44_add_69263[10:0] ^ p44_add_69263[19:9], p44_add_69263[20:12] ^ p44_add_69263[31:23] ^ p44_add_69263[8:0], p44_add_69263[11:2] ^ p44_add_69263[22:13] ^ p44_add_69263[31:22]} + (p45_and_69354_comb ^ p44_add_69263 & p44_add_69126 ^ p44_and_69258);
  assign p45_add_69336_comb = {p45_add_69314_comb[5:0] ^ p45_add_69314_comb[10:5] ^ p45_add_69314_comb[24:19], p45_add_69314_comb[31:27] ^ p45_add_69314_comb[4:0] ^ p45_add_69314_comb[18:14], p45_add_69314_comb[26:13] ^ p45_add_69314_comb[31:18] ^ p45_add_69314_comb[13:0], p45_add_69314_comb[12:6] ^ p45_add_69314_comb[17:11] ^ p45_add_69314_comb[31:25]} + (p45_add_69314_comb & p44_add_69220 ^ ~(p45_add_69314_comb | ~p44_add_69099));
  assign p45_not_69337_comb = ~p44_add_69220;
  assign p45_add_69359_comb = p45_add_69313_comb + p45_add_69358_comb;

  // Registers for pipe stage 45:
  reg [31:0] p45_add_69099;
  reg [31:0] p45_add_69314;
  reg [31:0] p45_add_69336;
  reg [31:0] p45_add_69127;
  reg [31:0] p45_add_69126;
  reg [31:0] p45_not_69337;
  reg [31:0] p45_concat_68872;
  reg [31:0] p45_add_69149;
  reg [31:0] p45_add_69263;
  reg [31:0] p45_add_69264;
  reg [31:0] p45_and_69354;
  reg [31:0] p45_add_69359;
  reg [31:0] p45_concat_68877;
  reg [31:0] p45_concat_68743;
  reg [3:0] p45_xor_68897;
  reg [31:0] p45_concat_69021;
  reg [31:0] p45_add_68761;
  reg [31:0] p45_add_68894;
  reg [31:0] p45_add_68540;
  reg [31:0] p45_add_68702;
  reg [31:0] p45_add_68522;
  reg [31:0] p45_add_68121;
  reg [31:0] p45_add_67611;
  always_ff @ (posedge clk) begin
    p45_add_69099 <= p44_add_69099;
    p45_add_69314 <= p45_add_69314_comb;
    p45_add_69336 <= p45_add_69336_comb;
    p45_add_69127 <= p44_add_69127;
    p45_add_69126 <= p44_add_69126;
    p45_not_69337 <= p45_not_69337_comb;
    p45_concat_68872 <= p44_concat_68872;
    p45_add_69149 <= p44_add_69149;
    p45_add_69263 <= p44_add_69263;
    p45_add_69264 <= p44_add_69264;
    p45_and_69354 <= p45_and_69354_comb;
    p45_add_69359 <= p45_add_69359_comb;
    p45_concat_68877 <= p44_concat_68877;
    p45_concat_68743 <= p44_concat_68743;
    p45_xor_68897 <= p44_xor_68897;
    p45_concat_69021 <= p44_concat_69021;
    p45_add_68761 <= p44_add_68761;
    p45_add_68894 <= p44_add_68894;
    p45_add_68540 <= p44_add_68540;
    p45_add_68702 <= p44_add_68702;
    p45_add_68522 <= p44_add_68522;
    p45_add_68121 <= p44_add_68121;
    p45_add_67611 <= p44_add_67611;
  end

  // ===== Pipe stage 46:
  wire [31:0] p46_add_69407_comb;
  wire [31:0] p46_add_69408_comb;
  wire [31:0] p46_add_69409_comb;
  wire [31:0] p46_and_69448_comb;
  wire [31:0] p46_add_69452_comb;
  wire [31:0] p46_add_69453_comb;
  wire [31:0] p46_add_69430_comb;
  wire [31:0] p46_add_69431_comb;
  assign p46_add_69407_comb = p45_add_69336 + 32'h391c_0cb3;
  assign p46_add_69408_comb = p46_add_69407_comb + p45_add_69127;
  assign p46_add_69409_comb = p45_add_69126 + p46_add_69408_comb;
  assign p46_and_69448_comb = p45_add_69359 & p45_add_69263;
  assign p46_add_69452_comb = {p45_add_69359[1:0] ^ p45_add_69359[12:11] ^ p45_add_69359[21:20], p45_add_69359[31:21] ^ p45_add_69359[10:0] ^ p45_add_69359[19:9], p45_add_69359[20:12] ^ p45_add_69359[31:23] ^ p45_add_69359[8:0], p45_add_69359[11:2] ^ p45_add_69359[22:13] ^ p45_add_69359[31:22]} + (p46_and_69448_comb ^ p45_add_69359 & p45_add_69149 ^ p45_and_69354);
  assign p46_add_69453_comb = p46_add_69408_comb + p46_add_69452_comb;
  assign p46_add_69430_comb = {p46_add_69409_comb[5:0] ^ p46_add_69409_comb[10:5] ^ p46_add_69409_comb[24:19], p46_add_69409_comb[31:27] ^ p46_add_69409_comb[4:0] ^ p46_add_69409_comb[18:14], p46_add_69409_comb[26:13] ^ p46_add_69409_comb[31:18] ^ p46_add_69409_comb[13:0], p46_add_69409_comb[12:6] ^ p46_add_69409_comb[17:11] ^ p46_add_69409_comb[31:25]} + p45_add_69099;
  assign p46_add_69431_comb = (p46_add_69409_comb & p45_add_69314 ^ ~(p46_add_69409_comb | p45_not_69337)) + p45_concat_68872;

  // Registers for pipe stage 46:
  reg [31:0] p46_add_69314;
  reg [31:0] p46_add_69409;
  reg [31:0] p46_add_69149;
  reg [31:0] p46_add_69263;
  reg [31:0] p46_add_69264;
  reg [31:0] p46_add_69359;
  reg [31:0] p46_and_69448;
  reg [31:0] p46_add_69453;
  reg [31:0] p46_concat_68877;
  reg [31:0] p46_concat_68743;
  reg [3:0] p46_xor_68897;
  reg [31:0] p46_concat_69021;
  reg [31:0] p46_add_68761;
  reg [31:0] p46_add_68894;
  reg [31:0] p46_add_68540;
  reg [31:0] p46_add_68702;
  reg [31:0] p46_add_68522;
  reg [31:0] p46_add_69430;
  reg [31:0] p46_add_69431;
  reg [31:0] p46_add_68121;
  reg [31:0] p46_add_67611;
  always_ff @ (posedge clk) begin
    p46_add_69314 <= p45_add_69314;
    p46_add_69409 <= p46_add_69409_comb;
    p46_add_69149 <= p45_add_69149;
    p46_add_69263 <= p45_add_69263;
    p46_add_69264 <= p45_add_69264;
    p46_add_69359 <= p45_add_69359;
    p46_and_69448 <= p46_and_69448_comb;
    p46_add_69453 <= p46_add_69453_comb;
    p46_concat_68877 <= p45_concat_68877;
    p46_concat_68743 <= p45_concat_68743;
    p46_xor_68897 <= p45_xor_68897;
    p46_concat_69021 <= p45_concat_69021;
    p46_add_68761 <= p45_add_68761;
    p46_add_68894 <= p45_add_68894;
    p46_add_68540 <= p45_add_68540;
    p46_add_68702 <= p45_add_68702;
    p46_add_68522 <= p45_add_68522;
    p46_add_69430 <= p46_add_69430_comb;
    p46_add_69431 <= p46_add_69431_comb;
    p46_add_68121 <= p45_add_68121;
    p46_add_67611 <= p45_add_67611;
  end

  // ===== Pipe stage 47:
  wire [31:0] p47_add_69496_comb;
  wire [31:0] p47_add_69497_comb;
  wire [31:0] p47_and_69539_comb;
  wire [31:0] p47_add_69543_comb;
  wire [31:0] p47_add_69519_comb;
  wire [31:0] p47_add_69522_comb;
  wire [31:0] p47_add_69544_comb;
  wire [31:0] p47_add_69545_comb;
  wire [31:0] p47_add_69521_comb;
  assign p47_add_69496_comb = p46_add_69430 + p46_add_69431;
  assign p47_add_69497_comb = p46_add_69149 + p47_add_69496_comb;
  assign p47_and_69539_comb = p46_add_69453 & p46_add_69359;
  assign p47_add_69543_comb = {p46_add_69453[1:0] ^ p46_add_69453[12:11] ^ p46_add_69453[21:20], p46_add_69453[31:21] ^ p46_add_69453[10:0] ^ p46_add_69453[19:9], p46_add_69453[20:12] ^ p46_add_69453[31:23] ^ p46_add_69453[8:0], p46_add_69453[11:2] ^ p46_add_69453[22:13] ^ p46_add_69453[31:22]} + (p47_and_69539_comb ^ p46_add_69453 & p46_add_69263 ^ p46_and_69448);
  assign p47_add_69519_comb = {p47_add_69497_comb[5:0] ^ p47_add_69497_comb[10:5] ^ p47_add_69497_comb[24:19], p47_add_69497_comb[31:27] ^ p47_add_69497_comb[4:0] ^ p47_add_69497_comb[18:14], p47_add_69497_comb[26:13] ^ p47_add_69497_comb[31:18] ^ p47_add_69497_comb[13:0], p47_add_69497_comb[12:6] ^ p47_add_69497_comb[17:11] ^ p47_add_69497_comb[31:25]} + (p47_add_69497_comb & p46_add_69409 ^ ~(p47_add_69497_comb | ~p46_add_69314));
  assign p47_add_69522_comb = p46_add_69314 + p46_add_68522;
  assign p47_add_69544_comb = p47_add_69496_comb + p47_add_69543_comb;
  assign p47_add_69545_comb = p47_add_69497_comb + p46_add_68540;
  assign p47_add_69521_comb = p47_add_69519_comb + 32'h5b9c_ca4f;

  // Registers for pipe stage 47:
  reg [31:0] p47_add_69409;
  reg [31:0] p47_add_69497;
  reg [31:0] p47_add_69263;
  reg [31:0] p47_add_69264;
  reg [31:0] p47_add_69359;
  reg [31:0] p47_add_69522;
  reg [31:0] p47_add_69453;
  reg [31:0] p47_and_69539;
  reg [31:0] p47_add_69544;
  reg [31:0] p47_add_69545;
  reg [31:0] p47_concat_68877;
  reg [31:0] p47_concat_68743;
  reg [3:0] p47_xor_68897;
  reg [31:0] p47_concat_69021;
  reg [31:0] p47_add_69521;
  reg [31:0] p47_add_68761;
  reg [31:0] p47_add_68894;
  reg [31:0] p47_add_68702;
  reg [31:0] p47_add_68522;
  reg [31:0] p47_add_68121;
  reg [31:0] p47_add_67611;
  always_ff @ (posedge clk) begin
    p47_add_69409 <= p46_add_69409;
    p47_add_69497 <= p47_add_69497_comb;
    p47_add_69263 <= p46_add_69263;
    p47_add_69264 <= p46_add_69264;
    p47_add_69359 <= p46_add_69359;
    p47_add_69522 <= p47_add_69522_comb;
    p47_add_69453 <= p46_add_69453;
    p47_and_69539 <= p47_and_69539_comb;
    p47_add_69544 <= p47_add_69544_comb;
    p47_add_69545 <= p47_add_69545_comb;
    p47_concat_68877 <= p46_concat_68877;
    p47_concat_68743 <= p46_concat_68743;
    p47_xor_68897 <= p46_xor_68897;
    p47_concat_69021 <= p46_concat_69021;
    p47_add_69521 <= p47_add_69521_comb;
    p47_add_68761 <= p46_add_68761;
    p47_add_68894 <= p46_add_68894;
    p47_add_68702 <= p46_add_68702;
    p47_add_68522 <= p46_add_68522;
    p47_add_68121 <= p46_add_68121;
    p47_add_67611 <= p46_add_67611;
  end

  // ===== Pipe stage 48:
  wire [31:0] p48_add_69588_comb;
  wire [31:0] p48_add_69589_comb;
  wire [31:0] p48_and_69631_comb;
  wire [31:0] p48_add_69635_comb;
  wire [31:0] p48_add_69611_comb;
  wire [31:0] p48_not_69614_comb;
  wire [31:0] p48_add_69636_comb;
  wire [31:0] p48_add_69613_comb;
  assign p48_add_69588_comb = p47_add_69521 + p47_add_69264;
  assign p48_add_69589_comb = p47_add_69263 + p48_add_69588_comb;
  assign p48_and_69631_comb = p47_add_69544 & p47_add_69453;
  assign p48_add_69635_comb = {p47_add_69544[1:0] ^ p47_add_69544[12:11] ^ p47_add_69544[21:20], p47_add_69544[31:21] ^ p47_add_69544[10:0] ^ p47_add_69544[19:9], p47_add_69544[20:12] ^ p47_add_69544[31:23] ^ p47_add_69544[8:0], p47_add_69544[11:2] ^ p47_add_69544[22:13] ^ p47_add_69544[31:22]} + (p48_and_69631_comb ^ p47_add_69544 & p47_add_69359 ^ p47_and_69539);
  assign p48_add_69611_comb = {p48_add_69589_comb[5:0] ^ p48_add_69589_comb[10:5] ^ p48_add_69589_comb[24:19], p48_add_69589_comb[31:27] ^ p48_add_69589_comb[4:0] ^ p48_add_69589_comb[18:14], p48_add_69589_comb[26:13] ^ p48_add_69589_comb[31:18] ^ p48_add_69589_comb[13:0], p48_add_69589_comb[12:6] ^ p48_add_69589_comb[17:11] ^ p48_add_69589_comb[31:25]} + (p48_add_69589_comb & p47_add_69497 ^ ~(p48_add_69589_comb | ~p47_add_69409));
  assign p48_not_69614_comb = ~p47_add_69497;
  assign p48_add_69636_comb = p48_add_69588_comb + p48_add_69635_comb;
  assign p48_add_69613_comb = p48_add_69611_comb + 32'h682e_6ff3;

  // Registers for pipe stage 48:
  reg [31:0] p48_add_69409;
  reg [31:0] p48_add_69589;
  reg [31:0] p48_add_69359;
  reg [31:0] p48_add_69522;
  reg [31:0] p48_not_69614;
  reg [31:0] p48_add_69453;
  reg [31:0] p48_add_69544;
  reg [31:0] p48_and_69631;
  reg [31:0] p48_add_69636;
  reg [31:0] p48_add_69545;
  reg [31:0] p48_concat_68877;
  reg [31:0] p48_concat_68743;
  reg [3:0] p48_xor_68897;
  reg [31:0] p48_concat_69021;
  reg [31:0] p48_add_69613;
  reg [31:0] p48_add_68761;
  reg [31:0] p48_add_68894;
  reg [31:0] p48_add_68702;
  reg [31:0] p48_add_68522;
  reg [31:0] p48_add_68121;
  reg [31:0] p48_add_67611;
  always_ff @ (posedge clk) begin
    p48_add_69409 <= p47_add_69409;
    p48_add_69589 <= p48_add_69589_comb;
    p48_add_69359 <= p47_add_69359;
    p48_add_69522 <= p47_add_69522;
    p48_not_69614 <= p48_not_69614_comb;
    p48_add_69453 <= p47_add_69453;
    p48_add_69544 <= p47_add_69544;
    p48_and_69631 <= p48_and_69631_comb;
    p48_add_69636 <= p48_add_69636_comb;
    p48_add_69545 <= p47_add_69545;
    p48_concat_68877 <= p47_concat_68877;
    p48_concat_68743 <= p47_concat_68743;
    p48_xor_68897 <= p47_xor_68897;
    p48_concat_69021 <= p47_concat_69021;
    p48_add_69613 <= p48_add_69613_comb;
    p48_add_68761 <= p47_add_68761;
    p48_add_68894 <= p47_add_68894;
    p48_add_68702 <= p47_add_68702;
    p48_add_68522 <= p47_add_68522;
    p48_add_68121 <= p47_add_68121;
    p48_add_67611 <= p47_add_67611;
  end

  // ===== Pipe stage 49:
  wire [31:0] p49_add_69679_comb;
  wire [31:0] p49_add_69680_comb;
  wire [31:0] p49_and_69725_comb;
  wire [30:0] p49_add_69701_comb;
  wire [31:0] p49_add_69729_comb;
  wire [31:0] p49_add_69706_comb;
  wire [31:0] p49_add_69707_comb;
  wire [31:0] p49_add_69730_comb;
  wire [31:0] p49_add_69708_comb;
  assign p49_add_69679_comb = p48_add_69613 + p48_add_69522;
  assign p49_add_69680_comb = p48_add_69359 + p49_add_69679_comb;
  assign p49_and_69725_comb = p48_add_69636 & p48_add_69544;
  assign p49_add_69701_comb = p48_add_68702[31:1] + 31'h3a47_c177;
  assign p49_add_69729_comb = {p48_add_69636[1:0] ^ p48_add_69636[12:11] ^ p48_add_69636[21:20], p48_add_69636[31:21] ^ p48_add_69636[10:0] ^ p48_add_69636[19:9], p48_add_69636[20:12] ^ p48_add_69636[31:23] ^ p48_add_69636[8:0], p48_add_69636[11:2] ^ p48_add_69636[22:13] ^ p48_add_69636[31:22]} + (p49_and_69725_comb ^ p48_add_69636 & p48_add_69453 ^ p48_and_69631);
  assign p49_add_69706_comb = {p49_add_69680_comb[5:0] ^ p49_add_69680_comb[10:5] ^ p49_add_69680_comb[24:19], p49_add_69680_comb[31:27] ^ p49_add_69680_comb[4:0] ^ p49_add_69680_comb[18:14], p49_add_69680_comb[26:13] ^ p49_add_69680_comb[31:18] ^ p49_add_69680_comb[13:0], p49_add_69680_comb[12:6] ^ p49_add_69680_comb[17:11] ^ p49_add_69680_comb[31:25]} + p48_add_69409;
  assign p49_add_69707_comb = (p49_add_69680_comb & p48_add_69589 ^ ~(p49_add_69680_comb | p48_not_69614)) + {p49_add_69701_comb, p48_add_68702[0]};
  assign p49_add_69730_comb = p49_add_69679_comb + p49_add_69729_comb;
  assign p49_add_69708_comb = p49_add_69706_comb + p49_add_69707_comb;

  // Registers for pipe stage 49:
  reg [31:0] p49_add_69589;
  reg [31:0] p49_add_69680;
  reg [31:0] p49_add_69453;
  reg [31:0] p49_add_69544;
  reg [31:0] p49_add_69636;
  reg [31:0] p49_add_69545;
  reg [31:0] p49_and_69725;
  reg [31:0] p49_concat_68877;
  reg [31:0] p49_add_69730;
  reg [31:0] p49_concat_68743;
  reg [3:0] p49_xor_68897;
  reg [31:0] p49_concat_69021;
  reg [31:0] p49_add_68761;
  reg [31:0] p49_add_68894;
  reg [31:0] p49_add_69708;
  reg [31:0] p49_add_68702;
  reg [31:0] p49_add_68522;
  reg [31:0] p49_add_68121;
  reg [31:0] p49_add_67611;
  always_ff @ (posedge clk) begin
    p49_add_69589 <= p48_add_69589;
    p49_add_69680 <= p49_add_69680_comb;
    p49_add_69453 <= p48_add_69453;
    p49_add_69544 <= p48_add_69544;
    p49_add_69636 <= p48_add_69636;
    p49_add_69545 <= p48_add_69545;
    p49_and_69725 <= p49_and_69725_comb;
    p49_concat_68877 <= p48_concat_68877;
    p49_add_69730 <= p49_add_69730_comb;
    p49_concat_68743 <= p48_concat_68743;
    p49_xor_68897 <= p48_xor_68897;
    p49_concat_69021 <= p48_concat_69021;
    p49_add_68761 <= p48_add_68761;
    p49_add_68894 <= p48_add_68894;
    p49_add_69708 <= p49_add_69708_comb;
    p49_add_68702 <= p48_add_68702;
    p49_add_68522 <= p48_add_68522;
    p49_add_68121 <= p48_add_68121;
    p49_add_67611 <= p48_add_67611;
  end

  // ===== Pipe stage 50:
  wire [31:0] p50_add_69769_comb;
  wire [31:0] p50_and_69811_comb;
  wire [31:0] p50_add_69791_comb;
  wire [31:0] p50_add_69793_comb;
  wire [31:0] p50_add_69815_comb;
  wire [31:0] p50_add_69794_comb;
  wire [31:0] p50_add_69816_comb;
  assign p50_add_69769_comb = p49_add_69453 + p49_add_69708;
  assign p50_and_69811_comb = p49_add_69730 & p49_add_69636;
  assign p50_add_69791_comb = {p50_add_69769_comb[5:0] ^ p50_add_69769_comb[10:5] ^ p50_add_69769_comb[24:19], p50_add_69769_comb[31:27] ^ p50_add_69769_comb[4:0] ^ p50_add_69769_comb[18:14], p50_add_69769_comb[26:13] ^ p50_add_69769_comb[31:18] ^ p50_add_69769_comb[13:0], p50_add_69769_comb[12:6] ^ p50_add_69769_comb[17:11] ^ p50_add_69769_comb[31:25]} + (p50_add_69769_comb & p49_add_69680 ^ ~(p50_add_69769_comb | ~p49_add_69589));
  assign p50_add_69793_comb = p50_add_69791_comb + 32'h78a5_636f;
  assign p50_add_69815_comb = {p49_add_69730[1:0] ^ p49_add_69730[12:11] ^ p49_add_69730[21:20], p49_add_69730[31:21] ^ p49_add_69730[10:0] ^ p49_add_69730[19:9], p49_add_69730[20:12] ^ p49_add_69730[31:23] ^ p49_add_69730[8:0], p49_add_69730[11:2] ^ p49_add_69730[22:13] ^ p49_add_69730[31:22]} + (p50_and_69811_comb ^ p49_add_69730 & p49_add_69544 ^ p49_and_69725);
  assign p50_add_69794_comb = p50_add_69793_comb + p49_add_69545;
  assign p50_add_69816_comb = p49_add_69708 + p50_add_69815_comb;

  // Registers for pipe stage 50:
  reg [31:0] p50_add_69589;
  reg [31:0] p50_add_69680;
  reg [31:0] p50_add_69544;
  reg [31:0] p50_add_69769;
  reg [31:0] p50_add_69636;
  reg [31:0] p50_add_69794;
  reg [31:0] p50_concat_68877;
  reg [31:0] p50_add_69730;
  reg [31:0] p50_and_69811;
  reg [31:0] p50_add_69816;
  reg [31:0] p50_concat_68743;
  reg [3:0] p50_xor_68897;
  reg [31:0] p50_concat_69021;
  reg [31:0] p50_add_68761;
  reg [31:0] p50_add_68894;
  reg [31:0] p50_add_68702;
  reg [31:0] p50_add_68522;
  reg [31:0] p50_add_68121;
  reg [31:0] p50_add_67611;
  always_ff @ (posedge clk) begin
    p50_add_69589 <= p49_add_69589;
    p50_add_69680 <= p49_add_69680;
    p50_add_69544 <= p49_add_69544;
    p50_add_69769 <= p50_add_69769_comb;
    p50_add_69636 <= p49_add_69636;
    p50_add_69794 <= p50_add_69794_comb;
    p50_concat_68877 <= p49_concat_68877;
    p50_add_69730 <= p49_add_69730;
    p50_and_69811 <= p50_and_69811_comb;
    p50_add_69816 <= p50_add_69816_comb;
    p50_concat_68743 <= p49_concat_68743;
    p50_xor_68897 <= p49_xor_68897;
    p50_concat_69021 <= p49_concat_69021;
    p50_add_68761 <= p49_add_68761;
    p50_add_68894 <= p49_add_68894;
    p50_add_68702 <= p49_add_68702;
    p50_add_68522 <= p49_add_68522;
    p50_add_68121 <= p49_add_68121;
    p50_add_67611 <= p49_add_67611;
  end

  // ===== Pipe stage 51:
  wire [31:0] p51_and_69897_comb;
  wire [31:0] p51_add_69855_comb;
  wire [31:0] p51_add_69901_comb;
  wire [31:0] p51_add_69902_comb;
  wire [31:0] p51_and_69919_comb;
  wire [31:0] p51_add_69877_comb;
  wire [31:0] p51_add_69878_comb;
  wire [31:0] p51_add_69879_comb;
  wire [31:0] p51_add_69923_comb;
  wire [31:0] p51_add_69892_comb;
  wire [31:0] p51_add_69924_comb;
  assign p51_and_69897_comb = p50_add_69816 & p50_add_69730;
  assign p51_add_69855_comb = p50_add_69544 + p50_add_69794;
  assign p51_add_69901_comb = {p50_add_69816[1:0] ^ p50_add_69816[12:11] ^ p50_add_69816[21:20], p50_add_69816[31:21] ^ p50_add_69816[10:0] ^ p50_add_69816[19:9], p50_add_69816[20:12] ^ p50_add_69816[31:23] ^ p50_add_69816[8:0], p50_add_69816[11:2] ^ p50_add_69816[22:13] ^ p50_add_69816[31:22]} + (p51_and_69897_comb ^ p50_add_69816 & p50_add_69636 ^ p50_and_69811);
  assign p51_add_69902_comb = p50_add_69794 + p51_add_69901_comb;
  assign p51_and_69919_comb = p51_add_69902_comb & p50_add_69816;
  assign p51_add_69877_comb = {p51_add_69855_comb[5:0] ^ p51_add_69855_comb[10:5] ^ p51_add_69855_comb[24:19], p51_add_69855_comb[31:27] ^ p51_add_69855_comb[4:0] ^ p51_add_69855_comb[18:14], p51_add_69855_comb[26:13] ^ p51_add_69855_comb[31:18] ^ p51_add_69855_comb[13:0], p51_add_69855_comb[12:6] ^ p51_add_69855_comb[17:11] ^ p51_add_69855_comb[31:25]} + p50_add_69589;
  assign p51_add_69878_comb = (p51_add_69855_comb & p50_add_69769 ^ ~(p51_add_69855_comb | ~p50_add_69680)) + p50_concat_68877;
  assign p51_add_69879_comb = p51_add_69877_comb + p51_add_69878_comb;
  assign p51_add_69923_comb = {p51_add_69902_comb[1:0] ^ p51_add_69902_comb[12:11] ^ p51_add_69902_comb[21:20], p51_add_69902_comb[31:21] ^ p51_add_69902_comb[10:0] ^ p51_add_69902_comb[19:9], p51_add_69902_comb[20:12] ^ p51_add_69902_comb[31:23] ^ p51_add_69902_comb[8:0], p51_add_69902_comb[11:2] ^ p51_add_69902_comb[22:13] ^ p51_add_69902_comb[31:22]} + (p51_and_69919_comb ^ p51_add_69902_comb & p50_add_69730 ^ p51_and_69897_comb);
  assign p51_add_69892_comb = p50_add_69636 + p51_add_69879_comb;
  assign p51_add_69924_comb = p51_add_69879_comb + p51_add_69923_comb;

  // Registers for pipe stage 51:
  reg [31:0] p51_add_69680;
  reg [31:0] p51_add_69769;
  reg [31:0] p51_add_69855;
  reg [31:0] p51_add_69730;
  reg [31:0] p51_add_69892;
  reg [31:0] p51_add_69816;
  reg [31:0] p51_concat_68743;
  reg [31:0] p51_add_69902;
  reg [31:0] p51_and_69919;
  reg [31:0] p51_add_69924;
  reg [3:0] p51_xor_68897;
  reg [31:0] p51_concat_69021;
  reg [31:0] p51_add_68761;
  reg [31:0] p51_add_68894;
  reg [31:0] p51_add_68702;
  reg [31:0] p51_add_68522;
  reg [31:0] p51_add_68121;
  reg [31:0] p51_add_67611;
  always_ff @ (posedge clk) begin
    p51_add_69680 <= p50_add_69680;
    p51_add_69769 <= p50_add_69769;
    p51_add_69855 <= p51_add_69855_comb;
    p51_add_69730 <= p50_add_69730;
    p51_add_69892 <= p51_add_69892_comb;
    p51_add_69816 <= p50_add_69816;
    p51_concat_68743 <= p50_concat_68743;
    p51_add_69902 <= p51_add_69902_comb;
    p51_and_69919 <= p51_and_69919_comb;
    p51_add_69924 <= p51_add_69924_comb;
    p51_xor_68897 <= p50_xor_68897;
    p51_concat_69021 <= p50_concat_69021;
    p51_add_68761 <= p50_add_68761;
    p51_add_68894 <= p50_add_68894;
    p51_add_68702 <= p50_add_68702;
    p51_add_68522 <= p50_add_68522;
    p51_add_68121 <= p50_add_68121;
    p51_add_67611 <= p50_add_67611;
  end

  // ===== Pipe stage 52:
  wire [31:0] p52_add_69982_comb;
  wire [31:0] p52_add_69983_comb;
  wire [31:0] p52_add_69984_comb;
  wire [12:0] p52_xor_70068_comb;
  wire [31:0] p52_add_69985_comb;
  wire [31:0] p52_and_70030_comb;
  wire [30:0] p52_add_70007_comb;
  wire [31:0] p52_add_70034_comb;
  wire [30:0] p52_add_70075_comb;
  wire [31:0] p52_not_70035_comb;
  wire [31:0] p52_add_70036_comb;
  wire [31:0] p52_add_70037_comb;
  wire [31:0] p52_concat_70077_comb;
  wire [31:0] p52_add_70078_comb;
  wire [31:0] p52_add_70055_comb;
  wire [31:0] p52_add_70056_comb;
  wire [31:0] p52_add_70024_comb;
  wire [31:0] p52_add_70025_comb;
  assign p52_add_69982_comb = {p51_add_69892[5:0] ^ p51_add_69892[10:5] ^ p51_add_69892[24:19], p51_add_69892[31:27] ^ p51_add_69892[4:0] ^ p51_add_69892[18:14], p51_add_69892[26:13] ^ p51_add_69892[31:18] ^ p51_add_69892[13:0], p51_add_69892[12:6] ^ p51_add_69892[17:11] ^ p51_add_69892[31:25]} + p51_add_69680;
  assign p52_add_69983_comb = (p51_add_69892 & p51_add_69855 ^ ~(p51_add_69892 | ~p51_add_69769)) + p51_concat_68743;
  assign p52_add_69984_comb = p52_add_69982_comb + p52_add_69983_comb;
  assign p52_xor_70068_comb = p51_add_68761[29:17] ^ p51_add_68761[31:19] ^ p51_add_68761[22:10];
  assign p52_add_69985_comb = p51_add_69730 + p52_add_69984_comb;
  assign p52_and_70030_comb = p51_add_69924 & p51_add_69902;
  assign p52_add_70007_comb = p51_add_68894[31:1] + 31'h485f_7ffd;
  assign p52_add_70034_comb = {p51_add_69924[1:0] ^ p51_add_69924[12:11] ^ p51_add_69924[21:20], p51_add_69924[31:21] ^ p51_add_69924[10:0] ^ p51_add_69924[19:9], p51_add_69924[20:12] ^ p51_add_69924[31:23] ^ p51_add_69924[8:0], p51_add_69924[11:2] ^ p51_add_69924[22:13] ^ p51_add_69924[31:22]} + (p52_and_70030_comb ^ p51_add_69924 & p51_add_69816 ^ p51_and_69919);
  assign p52_add_70075_comb = {p51_add_68761[16:7] ^ p51_add_68761[18:9], p51_add_68761[6:0] ^ p51_add_68761[8:2] ^ p51_add_68761[31:25], p51_add_68761[31:30] ^ p51_add_68761[1:0] ^ p51_add_68761[24:23], p52_xor_70068_comb[12:1]} + 31'h6338_bc79;
  assign p52_not_70035_comb = ~p51_add_69892;
  assign p52_add_70036_comb = p52_add_69984_comb + p52_add_70034_comb;
  assign p52_add_70037_comb = p51_add_69855 + p51_add_68761;
  assign p52_concat_70077_comb = {p52_add_70075_comb, p52_xor_70068_comb[0]};
  assign p52_add_70078_comb = p51_concat_69021 + p52_add_69985_comb;
  assign p52_add_70055_comb = p51_add_69892 + p51_add_68522;
  assign p52_add_70056_comb = {p51_add_68894[16:7] ^ p51_add_68894[18:9], p51_add_68894[6:0] ^ p51_add_68894[8:2] ^ p51_add_68894[31:25], p51_add_68894[31:30] ^ p51_add_68894[1:0] ^ p51_add_68894[24:23], p51_add_68894[29:17] ^ p51_add_68894[31:19] ^ p51_add_68894[22:10]} + 32'hbef9_a3f7;
  assign p52_add_70024_comb = {p52_add_69985_comb[5:0] ^ p52_add_69985_comb[10:5] ^ p52_add_69985_comb[24:19], p52_add_69985_comb[31:27] ^ p52_add_69985_comb[4:0] ^ p52_add_69985_comb[18:14], p52_add_69985_comb[26:13] ^ p52_add_69985_comb[31:18] ^ p52_add_69985_comb[13:0], p52_add_69985_comb[12:6] ^ p52_add_69985_comb[17:11] ^ p52_add_69985_comb[31:25]} + p51_add_69769;
  assign p52_add_70025_comb = (p52_add_69985_comb & p51_add_69892 ^ ~(p52_add_69985_comb | ~p51_add_69855)) + {p52_add_70007_comb, p51_add_68894[0]};

  // Registers for pipe stage 52:
  reg [31:0] p52_add_69816;
  reg [31:0] p52_add_69985;
  reg [31:0] p52_add_69902;
  reg [31:0] p52_add_69924;
  reg [31:0] p52_not_70035;
  reg [31:0] p52_and_70030;
  reg [31:0] p52_add_70036;
  reg [31:0] p52_add_70037;
  reg [3:0] p52_xor_68897;
  reg [31:0] p52_concat_70077;
  reg [31:0] p52_add_70078;
  reg [31:0] p52_add_70055;
  reg [31:0] p52_add_70056;
  reg [31:0] p52_add_70024;
  reg [31:0] p52_add_70025;
  reg [31:0] p52_add_68702;
  reg [31:0] p52_add_68121;
  reg [31:0] p52_add_67611;
  always_ff @ (posedge clk) begin
    p52_add_69816 <= p51_add_69816;
    p52_add_69985 <= p52_add_69985_comb;
    p52_add_69902 <= p51_add_69902;
    p52_add_69924 <= p51_add_69924;
    p52_not_70035 <= p52_not_70035_comb;
    p52_and_70030 <= p52_and_70030_comb;
    p52_add_70036 <= p52_add_70036_comb;
    p52_add_70037 <= p52_add_70037_comb;
    p52_xor_68897 <= p51_xor_68897;
    p52_concat_70077 <= p52_concat_70077_comb;
    p52_add_70078 <= p52_add_70078_comb;
    p52_add_70055 <= p52_add_70055_comb;
    p52_add_70056 <= p52_add_70056_comb;
    p52_add_70024 <= p52_add_70024_comb;
    p52_add_70025 <= p52_add_70025_comb;
    p52_add_68702 <= p51_add_68702;
    p52_add_68121 <= p51_add_68121;
    p52_add_67611 <= p51_add_67611;
  end

  // ===== Pipe stage 53:
  wire [31:0] p53_add_70115_comb;
  wire [31:0] p53_add_70116_comb;
  wire [31:0] p53_and_70153_comb;
  wire [31:0] p53_add_70160_comb;
  wire [31:0] p53_add_70155_comb;
  wire [31:0] p53_not_70162_comb;
  wire [31:0] p53_add_70161_comb;
  wire [31:0] p53_add_70159_comb;
  assign p53_add_70115_comb = p52_add_70024 + p52_add_70025;
  assign p53_add_70116_comb = p52_add_69816 + p53_add_70115_comb;
  assign p53_and_70153_comb = p52_add_70036 & p52_add_69924;
  assign p53_add_70160_comb = {p52_add_70036[1:0] ^ p52_add_70036[12:11] ^ p52_add_70036[21:20], p52_add_70036[31:21] ^ p52_add_70036[10:0] ^ p52_add_70036[19:9], p52_add_70036[20:12] ^ p52_add_70036[31:23] ^ p52_add_70036[8:0], p52_add_70036[11:2] ^ p52_add_70036[22:13] ^ p52_add_70036[31:22]} + (p53_and_70153_comb ^ p52_add_70036 & p52_add_69902 ^ p52_and_70030);
  assign p53_add_70155_comb = {p53_add_70116_comb[5:0] ^ p53_add_70116_comb[10:5] ^ p53_add_70116_comb[24:19], p53_add_70116_comb[31:27] ^ p53_add_70116_comb[4:0] ^ p53_add_70116_comb[18:14], p53_add_70116_comb[26:13] ^ p53_add_70116_comb[31:18] ^ p53_add_70116_comb[13:0], p53_add_70116_comb[12:6] ^ p53_add_70116_comb[17:11] ^ p53_add_70116_comb[31:25]} + (p53_add_70116_comb & p52_add_69985 ^ ~(p53_add_70116_comb | p52_not_70035));
  assign p53_not_70162_comb = ~p52_add_69985;
  assign p53_add_70161_comb = p53_add_70115_comb + p53_add_70160_comb;
  assign p53_add_70159_comb = p53_add_70155_comb + 32'ha450_6ceb;

  // Registers for pipe stage 53:
  reg [31:0] p53_add_69902;
  reg [31:0] p53_add_69924;
  reg [31:0] p53_add_70116;
  reg [31:0] p53_add_70036;
  reg [31:0] p53_add_70037;
  reg [31:0] p53_and_70153;
  reg [31:0] p53_not_70162;
  reg [3:0] p53_xor_68897;
  reg [31:0] p53_add_70161;
  reg [31:0] p53_concat_70077;
  reg [31:0] p53_add_70159;
  reg [31:0] p53_add_70078;
  reg [31:0] p53_add_70055;
  reg [31:0] p53_add_70056;
  reg [31:0] p53_add_68702;
  reg [31:0] p53_add_68121;
  reg [31:0] p53_add_67611;
  always_ff @ (posedge clk) begin
    p53_add_69902 <= p52_add_69902;
    p53_add_69924 <= p52_add_69924;
    p53_add_70116 <= p53_add_70116_comb;
    p53_add_70036 <= p52_add_70036;
    p53_add_70037 <= p52_add_70037;
    p53_and_70153 <= p53_and_70153_comb;
    p53_not_70162 <= p53_not_70162_comb;
    p53_xor_68897 <= p52_xor_68897;
    p53_add_70161 <= p53_add_70161_comb;
    p53_concat_70077 <= p52_concat_70077;
    p53_add_70159 <= p53_add_70159_comb;
    p53_add_70078 <= p52_add_70078;
    p53_add_70055 <= p52_add_70055;
    p53_add_70056 <= p52_add_70056;
    p53_add_68702 <= p52_add_68702;
    p53_add_68121 <= p52_add_68121;
    p53_add_67611 <= p52_add_67611;
  end

  // ===== Pipe stage 54:
  wire [31:0] p54_add_70197_comb;
  wire [31:0] p54_add_70198_comb;
  wire [31:0] p54_and_70235_comb;
  wire [31:0] p54_add_70251_comb;
  wire [31:0] p54_add_70252_comb;
  wire [31:0] p54_add_70253_comb;
  wire [31:0] p54_add_70254_comb;
  wire [31:0] p54_add_70255_comb;
  wire [31:0] p54_add_70256_comb;
  assign p54_add_70197_comb = p53_add_70159 + p53_add_70037;
  assign p54_add_70198_comb = p53_add_69902 + p54_add_70197_comb;
  assign p54_and_70235_comb = p53_add_70161 & p53_add_70036;
  assign p54_add_70251_comb = {p53_add_70161[1:0] ^ p53_add_70161[12:11] ^ p53_add_70161[21:20], p53_add_70161[31:21] ^ p53_add_70161[10:0] ^ p53_add_70161[19:9], p53_add_70161[20:12] ^ p53_add_70161[31:23] ^ p53_add_70161[8:0], p53_add_70161[11:2] ^ p53_add_70161[22:13] ^ p53_add_70161[31:22]} + (p54_and_70235_comb ^ p53_add_70161 & p53_add_69924 ^ p53_and_70153);
  assign p54_add_70252_comb = {p54_add_70198_comb[5:0] ^ p54_add_70198_comb[10:5] ^ p54_add_70198_comb[24:19], p54_add_70198_comb[31:27] ^ p54_add_70198_comb[4:0] ^ p54_add_70198_comb[18:14], p54_add_70198_comb[26:13] ^ p54_add_70198_comb[31:18] ^ p54_add_70198_comb[13:0], p54_add_70198_comb[12:6] ^ p54_add_70198_comb[17:11] ^ p54_add_70198_comb[31:25]} + {p53_add_68121[6:4] ^ p53_add_68121[17:15], p53_xor_68897, p53_add_68121[31:21] ^ p53_add_68121[10:0] ^ p53_add_68121[27:17], p53_add_68121[20:7] ^ p53_add_68121[31:18] ^ p53_add_68121[16:3]};
  assign p54_add_70253_comb = (p54_add_70198_comb & p53_add_70116 ^ ~(p54_add_70198_comb | p53_not_70162)) + p53_add_67611;
  assign p54_add_70254_comb = p54_add_70197_comb + p54_add_70251_comb;
  assign p54_add_70255_comb = p53_add_70055 + p54_add_70252_comb;
  assign p54_add_70256_comb = p54_add_70253_comb + p53_add_70056;

  // Registers for pipe stage 54:
  reg [31:0] p54_add_69924;
  reg [31:0] p54_add_70116;
  reg [31:0] p54_add_70036;
  reg [31:0] p54_add_70198;
  reg [31:0] p54_add_70161;
  reg [31:0] p54_and_70235;
  reg [31:0] p54_add_70254;
  reg [31:0] p54_concat_70077;
  reg [31:0] p54_add_70078;
  reg [31:0] p54_add_70255;
  reg [31:0] p54_add_70256;
  reg [31:0] p54_add_68702;
  reg [31:0] p54_add_68121;
  always_ff @ (posedge clk) begin
    p54_add_69924 <= p53_add_69924;
    p54_add_70116 <= p53_add_70116;
    p54_add_70036 <= p53_add_70036;
    p54_add_70198 <= p54_add_70198_comb;
    p54_add_70161 <= p53_add_70161;
    p54_and_70235 <= p54_and_70235_comb;
    p54_add_70254 <= p54_add_70254_comb;
    p54_concat_70077 <= p53_concat_70077;
    p54_add_70078 <= p53_add_70078;
    p54_add_70255 <= p54_add_70255_comb;
    p54_add_70256 <= p54_add_70256_comb;
    p54_add_68702 <= p53_add_68702;
    p54_add_68121 <= p53_add_68121;
  end

  // ===== Pipe stage 55:
  wire [31:0] p55_and_70300_comb;
  wire [31:0] p55_add_70295_comb;
  wire [31:0] p55_add_70302_comb;
  wire [31:0] p55_add_70318_comb;
  wire [31:0] p55_add_70325_comb;
  wire [30:0] p55_add_70344_comb;
  wire [30:0] p55_add_70346_comb;
  wire [29:0] p55_add_70349_comb;
  wire [31:0] p55_add_70328_comb;
  wire [31:0] p55_add_70329_comb;
  wire [31:0] p55_add_70348_comb;
  wire [31:0] p55_concat_70353_comb;
  wire [31:0] p55_concat_70354_comb;
  wire [31:0] p55_concat_70355_comb;
  wire [31:0] p55_add_70356_comb;
  wire [31:0] p55_add_70357_comb;
  wire [31:0] p55_add_70343_comb;
  wire [31:0] p55_add_70330_comb;
  wire [31:0] p55_add_70331_comb;
  assign p55_and_70300_comb = p54_add_70254 & p54_add_70161;
  assign p55_add_70295_comb = p54_add_70255 + p54_add_70256;
  assign p55_add_70302_comb = p54_add_69924 + p55_add_70295_comb;
  assign p55_add_70318_comb = {p54_add_70254[1:0] ^ p54_add_70254[12:11] ^ p54_add_70254[21:20], p54_add_70254[31:21] ^ p54_add_70254[10:0] ^ p54_add_70254[19:9], p54_add_70254[20:12] ^ p54_add_70254[31:23] ^ p54_add_70254[8:0], p54_add_70254[11:2] ^ p54_add_70254[22:13] ^ p54_add_70254[31:22]} + (p55_and_70300_comb ^ p54_add_70254 & p54_add_70036 ^ p54_and_70235);
  assign p55_add_70325_comb = p55_add_70295_comb + p55_add_70318_comb;
  assign p55_add_70344_comb = p54_add_70254[31:1] + 31'h1e37_79b9;
  assign p55_add_70346_comb = p54_add_70161[31:1] + 31'h52a7_fa9d;
  assign p55_add_70349_comb = p55_add_70302_comb[31:2] + 30'h26c1_5a23;
  assign p55_add_70328_comb = {p55_add_70302_comb[5:0] ^ p55_add_70302_comb[10:5] ^ p55_add_70302_comb[24:19], p55_add_70302_comb[31:27] ^ p55_add_70302_comb[4:0] ^ p55_add_70302_comb[18:14], p55_add_70302_comb[26:13] ^ p55_add_70302_comb[31:18] ^ p55_add_70302_comb[13:0], p55_add_70302_comb[12:6] ^ p55_add_70302_comb[17:11] ^ p55_add_70302_comb[31:25]} + p54_add_68121;
  assign p55_add_70329_comb = p54_concat_70077 + (p55_add_70302_comb & p54_add_70198 ^ ~(p55_add_70302_comb | ~p54_add_70116));
  assign p55_add_70348_comb = p54_add_70036 + 32'h510e_527f;
  assign p55_concat_70353_comb = {p55_add_70344_comb, p54_add_70254[0]};
  assign p55_concat_70354_comb = {p55_add_70346_comb, p54_add_70161[0]};
  assign p55_concat_70355_comb = {p55_add_70349_comb, p55_add_70302_comb[1:0]};
  assign p55_add_70356_comb = p54_add_70198 + 32'h1f83_d9ab;
  assign p55_add_70357_comb = p54_add_70116 + 32'h5be0_cd19;
  assign p55_add_70343_comb = (p55_add_70325_comb & p54_add_70254 ^ p55_add_70325_comb & p54_add_70161 ^ p55_and_70300_comb) + 32'h6a09_e667;
  assign p55_add_70330_comb = p55_add_70328_comb + p54_add_70078;
  assign p55_add_70331_comb = p55_add_70329_comb + p54_add_68702;

  // Registers for pipe stage 55:
  reg [31:0] p55_add_70325;
  reg [31:0] p55_add_70348;
  reg [31:0] p55_concat_70353;
  reg [31:0] p55_concat_70354;
  reg [31:0] p55_concat_70355;
  reg [31:0] p55_add_70356;
  reg [31:0] p55_add_70357;
  reg [31:0] p55_add_70343;
  reg [31:0] p55_add_70330;
  reg [31:0] p55_add_70331;
  always_ff @ (posedge clk) begin
    p55_add_70325 <= p55_add_70325_comb;
    p55_add_70348 <= p55_add_70348_comb;
    p55_concat_70353 <= p55_concat_70353_comb;
    p55_concat_70354 <= p55_concat_70354_comb;
    p55_concat_70355 <= p55_concat_70355_comb;
    p55_add_70356 <= p55_add_70356_comb;
    p55_add_70357 <= p55_add_70357_comb;
    p55_add_70343 <= p55_add_70343_comb;
    p55_add_70330 <= p55_add_70330_comb;
    p55_add_70331 <= p55_add_70331_comb;
  end

  // ===== Pipe stage 56:
  wire [31:0] p56_add_70395_comb;
  wire [31:0] p56_add_70396_comb;
  wire [31:0] p56_add_70398_comb;
  wire [31:0] p56_add_70399_comb;
  wire [31:0] p56_add_70400_comb;
  wire [255:0] p56_tuple_70401_comb;
  assign p56_add_70395_comb = p55_add_70330 + p55_add_70331;
  assign p56_add_70396_comb = {p55_add_70325[1:0] ^ p55_add_70325[12:11] ^ p55_add_70325[21:20], p55_add_70325[31:21] ^ p55_add_70325[10:0] ^ p55_add_70325[19:9], p55_add_70325[20:12] ^ p55_add_70325[31:23] ^ p55_add_70325[8:0], p55_add_70325[11:2] ^ p55_add_70325[22:13] ^ p55_add_70325[31:22]} + p56_add_70395_comb;
  assign p56_add_70398_comb = p56_add_70396_comb + p55_add_70343;
  assign p56_add_70399_comb = p55_add_70325 + 32'hbb67_ae85;
  assign p56_add_70400_comb = p56_add_70395_comb + p55_add_70348;
  assign p56_tuple_70401_comb = {p56_add_70398_comb, p56_add_70399_comb, p55_concat_70353, p55_concat_70354, p56_add_70400_comb, p55_concat_70355, p55_add_70356, p55_add_70357};

  // Registers for pipe stage 56:
  reg [255:0] p56_tuple_70401;
  always_ff @ (posedge clk) begin
    p56_tuple_70401 <= p56_tuple_70401_comb;
  end
  assign out = p56_tuple_70401;
endmodule
