module xls_test(
  input wire clk,
  input wire [2047:0] f,
  output wire [2047:0] out
);
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_11b (input reg [31:0] lhs, input reg [10:0] rhs);
    begin
      umul32b_32b_x_11b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_12b (input reg [31:0] lhs, input reg [11:0] rhs);
    begin
      umul32b_32b_x_12b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_10b (input reg [31:0] lhs, input reg [9:0] rhs);
    begin
      umul32b_32b_x_10b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_8b (input reg [31:0] lhs, input reg [7:0] rhs);
    begin
      umul32b_32b_x_8b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [31:0] f_unflattened[64];
  assign f_unflattened[0] = f[31:0];
  assign f_unflattened[1] = f[63:32];
  assign f_unflattened[2] = f[95:64];
  assign f_unflattened[3] = f[127:96];
  assign f_unflattened[4] = f[159:128];
  assign f_unflattened[5] = f[191:160];
  assign f_unflattened[6] = f[223:192];
  assign f_unflattened[7] = f[255:224];
  assign f_unflattened[8] = f[287:256];
  assign f_unflattened[9] = f[319:288];
  assign f_unflattened[10] = f[351:320];
  assign f_unflattened[11] = f[383:352];
  assign f_unflattened[12] = f[415:384];
  assign f_unflattened[13] = f[447:416];
  assign f_unflattened[14] = f[479:448];
  assign f_unflattened[15] = f[511:480];
  assign f_unflattened[16] = f[543:512];
  assign f_unflattened[17] = f[575:544];
  assign f_unflattened[18] = f[607:576];
  assign f_unflattened[19] = f[639:608];
  assign f_unflattened[20] = f[671:640];
  assign f_unflattened[21] = f[703:672];
  assign f_unflattened[22] = f[735:704];
  assign f_unflattened[23] = f[767:736];
  assign f_unflattened[24] = f[799:768];
  assign f_unflattened[25] = f[831:800];
  assign f_unflattened[26] = f[863:832];
  assign f_unflattened[27] = f[895:864];
  assign f_unflattened[28] = f[927:896];
  assign f_unflattened[29] = f[959:928];
  assign f_unflattened[30] = f[991:960];
  assign f_unflattened[31] = f[1023:992];
  assign f_unflattened[32] = f[1055:1024];
  assign f_unflattened[33] = f[1087:1056];
  assign f_unflattened[34] = f[1119:1088];
  assign f_unflattened[35] = f[1151:1120];
  assign f_unflattened[36] = f[1183:1152];
  assign f_unflattened[37] = f[1215:1184];
  assign f_unflattened[38] = f[1247:1216];
  assign f_unflattened[39] = f[1279:1248];
  assign f_unflattened[40] = f[1311:1280];
  assign f_unflattened[41] = f[1343:1312];
  assign f_unflattened[42] = f[1375:1344];
  assign f_unflattened[43] = f[1407:1376];
  assign f_unflattened[44] = f[1439:1408];
  assign f_unflattened[45] = f[1471:1440];
  assign f_unflattened[46] = f[1503:1472];
  assign f_unflattened[47] = f[1535:1504];
  assign f_unflattened[48] = f[1567:1536];
  assign f_unflattened[49] = f[1599:1568];
  assign f_unflattened[50] = f[1631:1600];
  assign f_unflattened[51] = f[1663:1632];
  assign f_unflattened[52] = f[1695:1664];
  assign f_unflattened[53] = f[1727:1696];
  assign f_unflattened[54] = f[1759:1728];
  assign f_unflattened[55] = f[1791:1760];
  assign f_unflattened[56] = f[1823:1792];
  assign f_unflattened[57] = f[1855:1824];
  assign f_unflattened[58] = f[1887:1856];
  assign f_unflattened[59] = f[1919:1888];
  assign f_unflattened[60] = f[1951:1920];
  assign f_unflattened[61] = f[1983:1952];
  assign f_unflattened[62] = f[2015:1984];
  assign f_unflattened[63] = f[2047:2016];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_f[64];
  always_ff @ (posedge clk) begin
    p0_f <= f_unflattened;
  end

  // ===== Pipe stage 1:
  wire [31:0] p1_array_index_32895_comb;
  wire [31:0] p1_array_index_32896_comb;
  wire [31:0] p1_array_index_32897_comb;
  wire [31:0] p1_array_index_32898_comb;
  wire [31:0] p1_array_index_32907_comb;
  wire [31:0] p1_array_index_32908_comb;
  wire [31:0] p1_array_index_32909_comb;
  wire [31:0] p1_array_index_32910_comb;
  wire [31:0] p1_array_index_32911_comb;
  wire [31:0] p1_array_index_32912_comb;
  wire [31:0] p1_array_index_32913_comb;
  wire [31:0] p1_array_index_32914_comb;
  wire [31:0] p1_array_index_32919_comb;
  wire [31:0] p1_array_index_32920_comb;
  wire [31:0] p1_array_index_32921_comb;
  wire [31:0] p1_array_index_32922_comb;
  wire [31:0] p1_array_index_32927_comb;
  wire [31:0] p1_array_index_32928_comb;
  wire [31:0] p1_array_index_32929_comb;
  wire [31:0] p1_array_index_32930_comb;
  wire [31:0] p1_array_index_32935_comb;
  wire [31:0] p1_array_index_32936_comb;
  wire [31:0] p1_array_index_32937_comb;
  wire [31:0] p1_array_index_32938_comb;
  wire [31:0] p1_array_index_32943_comb;
  wire [31:0] p1_array_index_32944_comb;
  wire [31:0] p1_array_index_32945_comb;
  wire [31:0] p1_array_index_32946_comb;
  wire [31:0] p1_array_index_32955_comb;
  wire [31:0] p1_array_index_32956_comb;
  wire [31:0] p1_array_index_32957_comb;
  wire [31:0] p1_array_index_32958_comb;
  wire [31:0] p1_array_index_32965_comb;
  wire [31:0] p1_array_index_32966_comb;
  wire [20:0] p1_bit_slice_32973_comb;
  wire [20:0] p1_bit_slice_32974_comb;
  wire [20:0] p1_bit_slice_32975_comb;
  wire [20:0] p1_bit_slice_32976_comb;
  wire [31:0] p1_array_index_32979_comb;
  wire [31:0] p1_array_index_32980_comb;
  wire [31:0] p1_array_index_32985_comb;
  wire [31:0] p1_array_index_32986_comb;
  wire [20:0] p1_bit_slice_32989_comb;
  wire [20:0] p1_bit_slice_32990_comb;
  wire [20:0] p1_bit_slice_32991_comb;
  wire [20:0] p1_bit_slice_32992_comb;
  wire [31:0] p1_array_index_32997_comb;
  wire [31:0] p1_array_index_32998_comb;
  wire [31:0] p1_array_index_32999_comb;
  wire [31:0] p1_array_index_33000_comb;
  wire [31:0] p1_array_index_33001_comb;
  wire [31:0] p1_array_index_33002_comb;
  wire [20:0] p1_bit_slice_33011_comb;
  wire [20:0] p1_bit_slice_33012_comb;
  wire [20:0] p1_bit_slice_33013_comb;
  wire [20:0] p1_bit_slice_33014_comb;
  wire [31:0] p1_array_index_33017_comb;
  wire [31:0] p1_array_index_33018_comb;
  wire [31:0] p1_array_index_33021_comb;
  wire [31:0] p1_array_index_33022_comb;
  wire [20:0] p1_bit_slice_33029_comb;
  wire [20:0] p1_bit_slice_33030_comb;
  wire [20:0] p1_bit_slice_33033_comb;
  wire [20:0] p1_bit_slice_33034_comb;
  assign p1_array_index_32895_comb = p0_f[6'h09];
  assign p1_array_index_32896_comb = p0_f[6'h0f];
  assign p1_array_index_32897_comb = p0_f[6'h39];
  assign p1_array_index_32898_comb = p0_f[6'h3f];
  assign p1_array_index_32907_comb = p0_f[6'h29];
  assign p1_array_index_32908_comb = p0_f[6'h2f];
  assign p1_array_index_32909_comb = p0_f[6'h19];
  assign p1_array_index_32910_comb = p0_f[6'h1f];
  assign p1_array_index_32911_comb = p0_f[6'h0d];
  assign p1_array_index_32912_comb = p0_f[6'h0b];
  assign p1_array_index_32913_comb = p0_f[6'h3d];
  assign p1_array_index_32914_comb = p0_f[6'h3b];
  assign p1_array_index_32919_comb = p0_f[6'h2d];
  assign p1_array_index_32920_comb = p0_f[6'h2b];
  assign p1_array_index_32921_comb = p0_f[6'h1d];
  assign p1_array_index_32922_comb = p0_f[6'h1b];
  assign p1_array_index_32927_comb = p0_f[6'h11];
  assign p1_array_index_32928_comb = p0_f[6'h17];
  assign p1_array_index_32929_comb = p0_f[6'h31];
  assign p1_array_index_32930_comb = p0_f[6'h37];
  assign p1_array_index_32935_comb = p0_f[6'h15];
  assign p1_array_index_32936_comb = p0_f[6'h13];
  assign p1_array_index_32937_comb = p0_f[6'h35];
  assign p1_array_index_32938_comb = p0_f[6'h33];
  assign p1_array_index_32943_comb = p0_f[6'h0a];
  assign p1_array_index_32944_comb = p0_f[6'h0e];
  assign p1_array_index_32945_comb = p0_f[6'h3a];
  assign p1_array_index_32946_comb = p0_f[6'h3e];
  assign p1_array_index_32955_comb = p0_f[6'h2a];
  assign p1_array_index_32956_comb = p0_f[6'h2e];
  assign p1_array_index_32957_comb = p0_f[6'h1a];
  assign p1_array_index_32958_comb = p0_f[6'h1e];
  assign p1_array_index_32965_comb = p0_f[6'h01];
  assign p1_array_index_32966_comb = p0_f[6'h07];
  assign p1_bit_slice_32973_comb = p0_f[6'h0c][20:0];
  assign p1_bit_slice_32974_comb = p0_f[6'h08][20:0];
  assign p1_bit_slice_32975_comb = p0_f[6'h3c][20:0];
  assign p1_bit_slice_32976_comb = p0_f[6'h38][20:0];
  assign p1_array_index_32979_comb = p0_f[6'h21];
  assign p1_array_index_32980_comb = p0_f[6'h27];
  assign p1_array_index_32985_comb = p0_f[6'h05];
  assign p1_array_index_32986_comb = p0_f[6'h03];
  assign p1_bit_slice_32989_comb = p0_f[6'h2c][20:0];
  assign p1_bit_slice_32990_comb = p0_f[6'h28][20:0];
  assign p1_bit_slice_32991_comb = p0_f[6'h1c][20:0];
  assign p1_bit_slice_32992_comb = p0_f[6'h18][20:0];
  assign p1_array_index_32997_comb = p0_f[6'h25];
  assign p1_array_index_32998_comb = p0_f[6'h23];
  assign p1_array_index_32999_comb = p0_f[6'h12];
  assign p1_array_index_33000_comb = p0_f[6'h16];
  assign p1_array_index_33001_comb = p0_f[6'h32];
  assign p1_array_index_33002_comb = p0_f[6'h36];
  assign p1_bit_slice_33011_comb = p0_f[6'h14][20:0];
  assign p1_bit_slice_33012_comb = p0_f[6'h10][20:0];
  assign p1_bit_slice_33013_comb = p0_f[6'h34][20:0];
  assign p1_bit_slice_33014_comb = p0_f[6'h30][20:0];
  assign p1_array_index_33017_comb = p0_f[6'h02];
  assign p1_array_index_33018_comb = p0_f[6'h06];
  assign p1_array_index_33021_comb = p0_f[6'h22];
  assign p1_array_index_33022_comb = p0_f[6'h26];
  assign p1_bit_slice_33029_comb = p0_f[6'h04][20:0];
  assign p1_bit_slice_33030_comb = p0_f[6'h00][20:0];
  assign p1_bit_slice_33033_comb = p0_f[6'h24][20:0];
  assign p1_bit_slice_33034_comb = p0_f[6'h20][20:0];

  // Registers for pipe stage 1:
  reg [31:0] p1_array_index_32895;
  reg [31:0] p1_array_index_32896;
  reg [31:0] p1_array_index_32897;
  reg [31:0] p1_array_index_32898;
  reg [31:0] p1_array_index_32907;
  reg [31:0] p1_array_index_32908;
  reg [31:0] p1_array_index_32909;
  reg [31:0] p1_array_index_32910;
  reg [31:0] p1_array_index_32911;
  reg [31:0] p1_array_index_32912;
  reg [31:0] p1_array_index_32913;
  reg [31:0] p1_array_index_32914;
  reg [31:0] p1_array_index_32919;
  reg [31:0] p1_array_index_32920;
  reg [31:0] p1_array_index_32921;
  reg [31:0] p1_array_index_32922;
  reg [31:0] p1_array_index_32927;
  reg [31:0] p1_array_index_32928;
  reg [31:0] p1_array_index_32929;
  reg [31:0] p1_array_index_32930;
  reg [31:0] p1_array_index_32935;
  reg [31:0] p1_array_index_32936;
  reg [31:0] p1_array_index_32937;
  reg [31:0] p1_array_index_32938;
  reg [31:0] p1_array_index_32943;
  reg [31:0] p1_array_index_32944;
  reg [31:0] p1_array_index_32945;
  reg [31:0] p1_array_index_32946;
  reg [31:0] p1_array_index_32955;
  reg [31:0] p1_array_index_32956;
  reg [31:0] p1_array_index_32957;
  reg [31:0] p1_array_index_32958;
  reg [31:0] p1_array_index_32965;
  reg [31:0] p1_array_index_32966;
  reg [20:0] p1_bit_slice_32973;
  reg [20:0] p1_bit_slice_32974;
  reg [20:0] p1_bit_slice_32975;
  reg [20:0] p1_bit_slice_32976;
  reg [31:0] p1_array_index_32979;
  reg [31:0] p1_array_index_32980;
  reg [31:0] p1_array_index_32985;
  reg [31:0] p1_array_index_32986;
  reg [20:0] p1_bit_slice_32989;
  reg [20:0] p1_bit_slice_32990;
  reg [20:0] p1_bit_slice_32991;
  reg [20:0] p1_bit_slice_32992;
  reg [31:0] p1_array_index_32997;
  reg [31:0] p1_array_index_32998;
  reg [31:0] p1_array_index_32999;
  reg [31:0] p1_array_index_33000;
  reg [31:0] p1_array_index_33001;
  reg [31:0] p1_array_index_33002;
  reg [20:0] p1_bit_slice_33011;
  reg [20:0] p1_bit_slice_33012;
  reg [20:0] p1_bit_slice_33013;
  reg [20:0] p1_bit_slice_33014;
  reg [31:0] p1_array_index_33017;
  reg [31:0] p1_array_index_33018;
  reg [31:0] p1_array_index_33021;
  reg [31:0] p1_array_index_33022;
  reg [20:0] p1_bit_slice_33029;
  reg [20:0] p1_bit_slice_33030;
  reg [20:0] p1_bit_slice_33033;
  reg [20:0] p1_bit_slice_33034;
  always_ff @ (posedge clk) begin
    p1_array_index_32895 <= p1_array_index_32895_comb;
    p1_array_index_32896 <= p1_array_index_32896_comb;
    p1_array_index_32897 <= p1_array_index_32897_comb;
    p1_array_index_32898 <= p1_array_index_32898_comb;
    p1_array_index_32907 <= p1_array_index_32907_comb;
    p1_array_index_32908 <= p1_array_index_32908_comb;
    p1_array_index_32909 <= p1_array_index_32909_comb;
    p1_array_index_32910 <= p1_array_index_32910_comb;
    p1_array_index_32911 <= p1_array_index_32911_comb;
    p1_array_index_32912 <= p1_array_index_32912_comb;
    p1_array_index_32913 <= p1_array_index_32913_comb;
    p1_array_index_32914 <= p1_array_index_32914_comb;
    p1_array_index_32919 <= p1_array_index_32919_comb;
    p1_array_index_32920 <= p1_array_index_32920_comb;
    p1_array_index_32921 <= p1_array_index_32921_comb;
    p1_array_index_32922 <= p1_array_index_32922_comb;
    p1_array_index_32927 <= p1_array_index_32927_comb;
    p1_array_index_32928 <= p1_array_index_32928_comb;
    p1_array_index_32929 <= p1_array_index_32929_comb;
    p1_array_index_32930 <= p1_array_index_32930_comb;
    p1_array_index_32935 <= p1_array_index_32935_comb;
    p1_array_index_32936 <= p1_array_index_32936_comb;
    p1_array_index_32937 <= p1_array_index_32937_comb;
    p1_array_index_32938 <= p1_array_index_32938_comb;
    p1_array_index_32943 <= p1_array_index_32943_comb;
    p1_array_index_32944 <= p1_array_index_32944_comb;
    p1_array_index_32945 <= p1_array_index_32945_comb;
    p1_array_index_32946 <= p1_array_index_32946_comb;
    p1_array_index_32955 <= p1_array_index_32955_comb;
    p1_array_index_32956 <= p1_array_index_32956_comb;
    p1_array_index_32957 <= p1_array_index_32957_comb;
    p1_array_index_32958 <= p1_array_index_32958_comb;
    p1_array_index_32965 <= p1_array_index_32965_comb;
    p1_array_index_32966 <= p1_array_index_32966_comb;
    p1_bit_slice_32973 <= p1_bit_slice_32973_comb;
    p1_bit_slice_32974 <= p1_bit_slice_32974_comb;
    p1_bit_slice_32975 <= p1_bit_slice_32975_comb;
    p1_bit_slice_32976 <= p1_bit_slice_32976_comb;
    p1_array_index_32979 <= p1_array_index_32979_comb;
    p1_array_index_32980 <= p1_array_index_32980_comb;
    p1_array_index_32985 <= p1_array_index_32985_comb;
    p1_array_index_32986 <= p1_array_index_32986_comb;
    p1_bit_slice_32989 <= p1_bit_slice_32989_comb;
    p1_bit_slice_32990 <= p1_bit_slice_32990_comb;
    p1_bit_slice_32991 <= p1_bit_slice_32991_comb;
    p1_bit_slice_32992 <= p1_bit_slice_32992_comb;
    p1_array_index_32997 <= p1_array_index_32997_comb;
    p1_array_index_32998 <= p1_array_index_32998_comb;
    p1_array_index_32999 <= p1_array_index_32999_comb;
    p1_array_index_33000 <= p1_array_index_33000_comb;
    p1_array_index_33001 <= p1_array_index_33001_comb;
    p1_array_index_33002 <= p1_array_index_33002_comb;
    p1_bit_slice_33011 <= p1_bit_slice_33011_comb;
    p1_bit_slice_33012 <= p1_bit_slice_33012_comb;
    p1_bit_slice_33013 <= p1_bit_slice_33013_comb;
    p1_bit_slice_33014 <= p1_bit_slice_33014_comb;
    p1_array_index_33017 <= p1_array_index_33017_comb;
    p1_array_index_33018 <= p1_array_index_33018_comb;
    p1_array_index_33021 <= p1_array_index_33021_comb;
    p1_array_index_33022 <= p1_array_index_33022_comb;
    p1_bit_slice_33029 <= p1_bit_slice_33029_comb;
    p1_bit_slice_33030 <= p1_bit_slice_33030_comb;
    p1_bit_slice_33033 <= p1_bit_slice_33033_comb;
    p1_bit_slice_33034 <= p1_bit_slice_33034_comb;
  end

  // ===== Pipe stage 2:
  wire [31:0] p2_umul_33253_comb;
  wire [31:0] p2_umul_33255_comb;
  wire [31:0] p2_umul_33269_comb;
  wire [31:0] p2_umul_33271_comb;
  wire [31:0] p2_umul_33285_comb;
  wire [31:0] p2_umul_33287_comb;
  wire [31:0] p2_add_33164_comb;
  wire [31:0] p2_add_33167_comb;
  wire [31:0] p2_add_33174_comb;
  wire [31:0] p2_add_33177_comb;
  wire [31:0] p2_add_33179_comb;
  wire [31:0] p2_add_33182_comb;
  wire [31:0] p2_add_33197_comb;
  wire [31:0] p2_add_33200_comb;
  wire [31:0] p2_add_33220_comb;
  wire [31:0] p2_add_33223_comb;
  wire [31:0] p2_add_33229_comb;
  wire [31:0] p2_add_33232_comb;
  wire [31:0] p2_add_33244_comb;
  wire [31:0] p2_add_33247_comb;
  wire [31:0] p2_add_33260_comb;
  wire [31:0] p2_add_33263_comb;
  wire [31:0] p2_add_33280_comb;
  wire [31:0] p2_add_33283_comb;
  wire [26:0] p2_bit_slice_33265_comb;
  wire [26:0] p2_bit_slice_33266_comb;
  wire [26:0] p2_bit_slice_33275_comb;
  wire [26:0] p2_bit_slice_33276_comb;
  wire [26:0] p2_bit_slice_33291_comb;
  wire [26:0] p2_bit_slice_33292_comb;
  wire [31:0] p2_umul_33169_comb;
  wire [31:0] p2_umul_33170_comb;
  wire [31:0] p2_umul_33171_comb;
  wire [31:0] p2_umul_33172_comb;
  wire [31:0] p2_umul_33185_comb;
  wire [31:0] p2_umul_33186_comb;
  wire [31:0] p2_umul_33187_comb;
  wire [31:0] p2_umul_33188_comb;
  wire [31:0] p2_umul_33189_comb;
  wire [31:0] p2_umul_33190_comb;
  wire [31:0] p2_umul_33193_comb;
  wire [31:0] p2_umul_33194_comb;
  wire [31:0] p2_umul_33203_comb;
  wire [31:0] p2_umul_33204_comb;
  wire [31:0] p2_umul_33205_comb;
  wire [31:0] p2_umul_33206_comb;
  wire [31:0] p2_umul_33207_comb;
  wire [31:0] p2_umul_33208_comb;
  wire [31:0] p2_umul_33211_comb;
  wire [31:0] p2_umul_33212_comb;
  wire [31:0] p2_umul_33215_comb;
  wire [31:0] p2_umul_33216_comb;
  wire [31:0] p2_umul_33217_comb;
  wire [31:0] p2_umul_33218_comb;
  wire [31:0] p2_umul_33225_comb;
  wire [31:0] p2_umul_33226_comb;
  wire [31:0] p2_umul_33227_comb;
  wire [31:0] p2_umul_33228_comb;
  wire [31:0] p2_umul_33235_comb;
  wire [31:0] p2_umul_33236_comb;
  wire [31:0] p2_umul_33239_comb;
  wire [31:0] p2_umul_33240_comb;
  wire [31:0] p2_umul_33249_comb;
  wire [31:0] p2_umul_33250_comb;
  wire [31:0] p2_umul_33251_comb;
  wire [31:0] p2_umul_33252_comb;
  wire [31:0] p2_umul_33254_comb;
  wire [31:0] p2_umul_33256_comb;
  wire [31:0] p2_umul_33267_comb;
  wire [31:0] p2_umul_33268_comb;
  wire [31:0] p2_umul_33270_comb;
  wire [31:0] p2_umul_33272_comb;
  wire [31:0] p2_umul_33277_comb;
  wire [31:0] p2_umul_33278_comb;
  wire [31:0] p2_umul_33286_comb;
  wire [31:0] p2_umul_33288_comb;
  wire [31:0] p2_umul_33293_comb;
  wire [31:0] p2_umul_33294_comb;
  assign p2_umul_33253_comb = umul32b_32b_x_11b(p1_array_index_32943, 11'h620);
  assign p2_umul_33255_comb = umul32b_32b_x_11b(p1_array_index_32945, 11'h620);
  assign p2_umul_33269_comb = umul32b_32b_x_11b(p1_array_index_32955, 11'h620);
  assign p2_umul_33271_comb = umul32b_32b_x_11b(p1_array_index_32957, 11'h620);
  assign p2_umul_33285_comb = umul32b_32b_x_11b(p1_array_index_32999, 11'h620);
  assign p2_umul_33287_comb = umul32b_32b_x_11b(p1_array_index_33001, 11'h620);
  assign p2_add_33164_comb = p1_array_index_32895 + p1_array_index_32896;
  assign p2_add_33167_comb = p1_array_index_32897 + p1_array_index_32898;
  assign p2_add_33174_comb = p1_array_index_32907 + p1_array_index_32908;
  assign p2_add_33177_comb = p1_array_index_32909 + p1_array_index_32910;
  assign p2_add_33179_comb = p1_array_index_32911 + p1_array_index_32912;
  assign p2_add_33182_comb = p1_array_index_32913 + p1_array_index_32914;
  assign p2_add_33197_comb = p1_array_index_32919 + p1_array_index_32920;
  assign p2_add_33200_comb = p1_array_index_32921 + p1_array_index_32922;
  assign p2_add_33220_comb = p1_array_index_32927 + p1_array_index_32928;
  assign p2_add_33223_comb = p1_array_index_32929 + p1_array_index_32930;
  assign p2_add_33229_comb = p1_array_index_32935 + p1_array_index_32936;
  assign p2_add_33232_comb = p1_array_index_32937 + p1_array_index_32938;
  assign p2_add_33244_comb = p1_array_index_32943 + p1_array_index_32944;
  assign p2_add_33247_comb = p1_array_index_32945 + p1_array_index_32946;
  assign p2_add_33260_comb = p1_array_index_32955 + p1_array_index_32956;
  assign p2_add_33263_comb = p1_array_index_32957 + p1_array_index_32958;
  assign p2_add_33280_comb = p1_array_index_32999 + p1_array_index_33000;
  assign p2_add_33283_comb = p1_array_index_33001 + p1_array_index_33002;
  assign p2_bit_slice_33265_comb = p2_umul_33253_comb[31:5];
  assign p2_bit_slice_33266_comb = p2_umul_33255_comb[31:5];
  assign p2_bit_slice_33275_comb = p2_umul_33269_comb[31:5];
  assign p2_bit_slice_33276_comb = p2_umul_33271_comb[31:5];
  assign p2_bit_slice_33291_comb = p2_umul_33285_comb[31:5];
  assign p2_bit_slice_33292_comb = p2_umul_33287_comb[31:5];
  assign p2_umul_33169_comb = umul32b_32b_x_12b(p1_array_index_32895, 12'h8e4);
  assign p2_umul_33170_comb = umul32b_32b_x_10b(p2_add_33164_comb, 10'h235);
  assign p2_umul_33171_comb = umul32b_32b_x_12b(p1_array_index_32897, 12'h8e4);
  assign p2_umul_33172_comb = umul32b_32b_x_10b(p2_add_33167_comb, 10'h235);
  assign p2_umul_33185_comb = umul32b_32b_x_12b(p1_array_index_32907, 12'h8e4);
  assign p2_umul_33186_comb = umul32b_32b_x_10b(p2_add_33174_comb, 10'h235);
  assign p2_umul_33187_comb = umul32b_32b_x_12b(p1_array_index_32909, 12'h8e4);
  assign p2_umul_33188_comb = umul32b_32b_x_10b(p2_add_33177_comb, 10'h235);
  assign p2_umul_33189_comb = umul32b_32b_x_12b(p2_add_33179_comb, 12'h968);
  assign p2_umul_33190_comb = umul32b_32b_x_12b(p1_array_index_32896, 12'hd4e);
  assign p2_umul_33193_comb = umul32b_32b_x_12b(p2_add_33182_comb, 12'h968);
  assign p2_umul_33194_comb = umul32b_32b_x_12b(p1_array_index_32898, 12'hd4e);
  assign p2_umul_33203_comb = umul32b_32b_x_10b(p1_array_index_32911, 10'h31f);
  assign p2_umul_33204_comb = umul32b_32b_x_12b(p1_array_index_32912, 12'hfb1);
  assign p2_umul_33205_comb = umul32b_32b_x_10b(p1_array_index_32913, 10'h31f);
  assign p2_umul_33206_comb = umul32b_32b_x_12b(p1_array_index_32914, 12'hfb1);
  assign p2_umul_33207_comb = umul32b_32b_x_12b(p2_add_33197_comb, 12'h968);
  assign p2_umul_33208_comb = umul32b_32b_x_12b(p1_array_index_32908, 12'hd4e);
  assign p2_umul_33211_comb = umul32b_32b_x_12b(p2_add_33200_comb, 12'h968);
  assign p2_umul_33212_comb = umul32b_32b_x_12b(p1_array_index_32910, 12'hd4e);
  assign p2_umul_33215_comb = umul32b_32b_x_10b(p1_array_index_32919, 10'h31f);
  assign p2_umul_33216_comb = umul32b_32b_x_12b(p1_array_index_32920, 12'hfb1);
  assign p2_umul_33217_comb = umul32b_32b_x_10b(p1_array_index_32921, 10'h31f);
  assign p2_umul_33218_comb = umul32b_32b_x_12b(p1_array_index_32922, 12'hfb1);
  assign p2_umul_33225_comb = umul32b_32b_x_12b(p1_array_index_32927, 12'h8e4);
  assign p2_umul_33226_comb = umul32b_32b_x_10b(p2_add_33220_comb, 10'h235);
  assign p2_umul_33227_comb = umul32b_32b_x_12b(p1_array_index_32929, 12'h8e4);
  assign p2_umul_33228_comb = umul32b_32b_x_10b(p2_add_33223_comb, 10'h235);
  assign p2_umul_33235_comb = umul32b_32b_x_12b(p2_add_33229_comb, 12'h968);
  assign p2_umul_33236_comb = umul32b_32b_x_12b(p1_array_index_32928, 12'hd4e);
  assign p2_umul_33239_comb = umul32b_32b_x_12b(p2_add_33232_comb, 12'h968);
  assign p2_umul_33240_comb = umul32b_32b_x_12b(p1_array_index_32930, 12'hd4e);
  assign p2_umul_33249_comb = umul32b_32b_x_10b(p1_array_index_32935, 10'h31f);
  assign p2_umul_33250_comb = umul32b_32b_x_12b(p1_array_index_32936, 12'hfb1);
  assign p2_umul_33251_comb = umul32b_32b_x_10b(p1_array_index_32937, 10'h31f);
  assign p2_umul_33252_comb = umul32b_32b_x_12b(p1_array_index_32938, 12'hfb1);
  assign p2_umul_33254_comb = umul32b_32b_x_11b(p2_add_33244_comb, 11'h454);
  assign p2_umul_33256_comb = umul32b_32b_x_11b(p2_add_33247_comb, 11'h454);
  assign p2_umul_33267_comb = umul32b_32b_x_12b(p1_array_index_32944, 12'hec8);
  assign p2_umul_33268_comb = umul32b_32b_x_12b(p1_array_index_32946, 12'hec8);
  assign p2_umul_33270_comb = umul32b_32b_x_11b(p2_add_33260_comb, 11'h454);
  assign p2_umul_33272_comb = umul32b_32b_x_11b(p2_add_33263_comb, 11'h454);
  assign p2_umul_33277_comb = umul32b_32b_x_12b(p1_array_index_32956, 12'hec8);
  assign p2_umul_33278_comb = umul32b_32b_x_12b(p1_array_index_32958, 12'hec8);
  assign p2_umul_33286_comb = umul32b_32b_x_11b(p2_add_33280_comb, 11'h454);
  assign p2_umul_33288_comb = umul32b_32b_x_11b(p2_add_33283_comb, 11'h454);
  assign p2_umul_33293_comb = umul32b_32b_x_12b(p1_array_index_33000, 12'hec8);
  assign p2_umul_33294_comb = umul32b_32b_x_12b(p1_array_index_33002, 12'hec8);

  // Registers for pipe stage 2:
  reg [26:0] p2_bit_slice_33265;
  reg [26:0] p2_bit_slice_33266;
  reg [31:0] p2_array_index_32965;
  reg [31:0] p2_array_index_32966;
  reg [20:0] p2_bit_slice_32973;
  reg [20:0] p2_bit_slice_32974;
  reg [20:0] p2_bit_slice_32975;
  reg [20:0] p2_bit_slice_32976;
  reg [31:0] p2_array_index_32979;
  reg [31:0] p2_array_index_32980;
  reg [26:0] p2_bit_slice_33275;
  reg [26:0] p2_bit_slice_33276;
  reg [31:0] p2_array_index_32985;
  reg [31:0] p2_array_index_32986;
  reg [20:0] p2_bit_slice_32989;
  reg [20:0] p2_bit_slice_32990;
  reg [20:0] p2_bit_slice_32991;
  reg [20:0] p2_bit_slice_32992;
  reg [31:0] p2_array_index_32997;
  reg [31:0] p2_array_index_32998;
  reg [26:0] p2_bit_slice_33291;
  reg [26:0] p2_bit_slice_33292;
  reg [20:0] p2_bit_slice_33011;
  reg [20:0] p2_bit_slice_33012;
  reg [20:0] p2_bit_slice_33013;
  reg [20:0] p2_bit_slice_33014;
  reg [31:0] p2_array_index_33017;
  reg [31:0] p2_array_index_33018;
  reg [31:0] p2_array_index_33021;
  reg [31:0] p2_array_index_33022;
  reg [20:0] p2_bit_slice_33029;
  reg [20:0] p2_bit_slice_33030;
  reg [20:0] p2_bit_slice_33033;
  reg [20:0] p2_bit_slice_33034;
  reg [31:0] p2_umul_33169;
  reg [31:0] p2_umul_33170;
  reg [31:0] p2_umul_33171;
  reg [31:0] p2_umul_33172;
  reg [31:0] p2_umul_33185;
  reg [31:0] p2_umul_33186;
  reg [31:0] p2_umul_33187;
  reg [31:0] p2_umul_33188;
  reg [31:0] p2_umul_33189;
  reg [31:0] p2_umul_33190;
  reg [31:0] p2_umul_33193;
  reg [31:0] p2_umul_33194;
  reg [31:0] p2_umul_33203;
  reg [31:0] p2_umul_33204;
  reg [31:0] p2_umul_33205;
  reg [31:0] p2_umul_33206;
  reg [31:0] p2_umul_33207;
  reg [31:0] p2_umul_33208;
  reg [31:0] p2_umul_33211;
  reg [31:0] p2_umul_33212;
  reg [31:0] p2_umul_33215;
  reg [31:0] p2_umul_33216;
  reg [31:0] p2_umul_33217;
  reg [31:0] p2_umul_33218;
  reg [31:0] p2_umul_33225;
  reg [31:0] p2_umul_33226;
  reg [31:0] p2_umul_33227;
  reg [31:0] p2_umul_33228;
  reg [31:0] p2_umul_33235;
  reg [31:0] p2_umul_33236;
  reg [31:0] p2_umul_33239;
  reg [31:0] p2_umul_33240;
  reg [31:0] p2_umul_33249;
  reg [31:0] p2_umul_33250;
  reg [31:0] p2_umul_33251;
  reg [31:0] p2_umul_33252;
  reg [31:0] p2_umul_33254;
  reg [31:0] p2_umul_33256;
  reg [31:0] p2_umul_33267;
  reg [31:0] p2_umul_33268;
  reg [31:0] p2_umul_33270;
  reg [31:0] p2_umul_33272;
  reg [31:0] p2_umul_33277;
  reg [31:0] p2_umul_33278;
  reg [31:0] p2_umul_33286;
  reg [31:0] p2_umul_33288;
  reg [31:0] p2_umul_33293;
  reg [31:0] p2_umul_33294;
  always_ff @ (posedge clk) begin
    p2_bit_slice_33265 <= p2_bit_slice_33265_comb;
    p2_bit_slice_33266 <= p2_bit_slice_33266_comb;
    p2_array_index_32965 <= p1_array_index_32965;
    p2_array_index_32966 <= p1_array_index_32966;
    p2_bit_slice_32973 <= p1_bit_slice_32973;
    p2_bit_slice_32974 <= p1_bit_slice_32974;
    p2_bit_slice_32975 <= p1_bit_slice_32975;
    p2_bit_slice_32976 <= p1_bit_slice_32976;
    p2_array_index_32979 <= p1_array_index_32979;
    p2_array_index_32980 <= p1_array_index_32980;
    p2_bit_slice_33275 <= p2_bit_slice_33275_comb;
    p2_bit_slice_33276 <= p2_bit_slice_33276_comb;
    p2_array_index_32985 <= p1_array_index_32985;
    p2_array_index_32986 <= p1_array_index_32986;
    p2_bit_slice_32989 <= p1_bit_slice_32989;
    p2_bit_slice_32990 <= p1_bit_slice_32990;
    p2_bit_slice_32991 <= p1_bit_slice_32991;
    p2_bit_slice_32992 <= p1_bit_slice_32992;
    p2_array_index_32997 <= p1_array_index_32997;
    p2_array_index_32998 <= p1_array_index_32998;
    p2_bit_slice_33291 <= p2_bit_slice_33291_comb;
    p2_bit_slice_33292 <= p2_bit_slice_33292_comb;
    p2_bit_slice_33011 <= p1_bit_slice_33011;
    p2_bit_slice_33012 <= p1_bit_slice_33012;
    p2_bit_slice_33013 <= p1_bit_slice_33013;
    p2_bit_slice_33014 <= p1_bit_slice_33014;
    p2_array_index_33017 <= p1_array_index_33017;
    p2_array_index_33018 <= p1_array_index_33018;
    p2_array_index_33021 <= p1_array_index_33021;
    p2_array_index_33022 <= p1_array_index_33022;
    p2_bit_slice_33029 <= p1_bit_slice_33029;
    p2_bit_slice_33030 <= p1_bit_slice_33030;
    p2_bit_slice_33033 <= p1_bit_slice_33033;
    p2_bit_slice_33034 <= p1_bit_slice_33034;
    p2_umul_33169 <= p2_umul_33169_comb;
    p2_umul_33170 <= p2_umul_33170_comb;
    p2_umul_33171 <= p2_umul_33171_comb;
    p2_umul_33172 <= p2_umul_33172_comb;
    p2_umul_33185 <= p2_umul_33185_comb;
    p2_umul_33186 <= p2_umul_33186_comb;
    p2_umul_33187 <= p2_umul_33187_comb;
    p2_umul_33188 <= p2_umul_33188_comb;
    p2_umul_33189 <= p2_umul_33189_comb;
    p2_umul_33190 <= p2_umul_33190_comb;
    p2_umul_33193 <= p2_umul_33193_comb;
    p2_umul_33194 <= p2_umul_33194_comb;
    p2_umul_33203 <= p2_umul_33203_comb;
    p2_umul_33204 <= p2_umul_33204_comb;
    p2_umul_33205 <= p2_umul_33205_comb;
    p2_umul_33206 <= p2_umul_33206_comb;
    p2_umul_33207 <= p2_umul_33207_comb;
    p2_umul_33208 <= p2_umul_33208_comb;
    p2_umul_33211 <= p2_umul_33211_comb;
    p2_umul_33212 <= p2_umul_33212_comb;
    p2_umul_33215 <= p2_umul_33215_comb;
    p2_umul_33216 <= p2_umul_33216_comb;
    p2_umul_33217 <= p2_umul_33217_comb;
    p2_umul_33218 <= p2_umul_33218_comb;
    p2_umul_33225 <= p2_umul_33225_comb;
    p2_umul_33226 <= p2_umul_33226_comb;
    p2_umul_33227 <= p2_umul_33227_comb;
    p2_umul_33228 <= p2_umul_33228_comb;
    p2_umul_33235 <= p2_umul_33235_comb;
    p2_umul_33236 <= p2_umul_33236_comb;
    p2_umul_33239 <= p2_umul_33239_comb;
    p2_umul_33240 <= p2_umul_33240_comb;
    p2_umul_33249 <= p2_umul_33249_comb;
    p2_umul_33250 <= p2_umul_33250_comb;
    p2_umul_33251 <= p2_umul_33251_comb;
    p2_umul_33252 <= p2_umul_33252_comb;
    p2_umul_33254 <= p2_umul_33254_comb;
    p2_umul_33256 <= p2_umul_33256_comb;
    p2_umul_33267 <= p2_umul_33267_comb;
    p2_umul_33268 <= p2_umul_33268_comb;
    p2_umul_33270 <= p2_umul_33270_comb;
    p2_umul_33272 <= p2_umul_33272_comb;
    p2_umul_33277 <= p2_umul_33277_comb;
    p2_umul_33278 <= p2_umul_33278_comb;
    p2_umul_33286 <= p2_umul_33286_comb;
    p2_umul_33288 <= p2_umul_33288_comb;
    p2_umul_33293 <= p2_umul_33293_comb;
    p2_umul_33294 <= p2_umul_33294_comb;
  end

  // ===== Pipe stage 3:
  wire [26:0] p3_add_33593_comb;
  wire [26:0] p3_add_33594_comb;
  wire [26:0] p3_add_33671_comb;
  wire [26:0] p3_add_33672_comb;
  wire [26:0] p3_add_33909_comb;
  wire [26:0] p3_add_33910_comb;
  wire [29:0] p3_add_33463_comb;
  wire [29:0] p3_add_33465_comb;
  wire [29:0] p3_add_33477_comb;
  wire [29:0] p3_add_33479_comb;
  wire [29:0] p3_add_33563_comb;
  wire [29:0] p3_add_33565_comb;
  wire [20:0] p3_add_33610_comb;
  wire [20:0] p3_add_33616_comb;
  wire [20:0] p3_add_33698_comb;
  wire [20:0] p3_add_33704_comb;
  wire [20:0] p3_add_33922_comb;
  wire [20:0] p3_add_33928_comb;
  wire [31:0] p3_concat_33473_comb;
  wire [31:0] p3_concat_33476_comb;
  wire [31:0] p3_concat_33491_comb;
  wire [31:0] p3_concat_33494_comb;
  wire [31:0] p3_concat_33573_comb;
  wire [31:0] p3_concat_33576_comb;
  wire [24:0] p3_add_33647_comb;
  wire [20:0] p3_add_33649_comb;
  wire [30:0] p3_add_33651_comb;
  wire [24:0] p3_add_33653_comb;
  wire [20:0] p3_add_33655_comb;
  wire [30:0] p3_add_33657_comb;
  wire [24:0] p3_add_33659_comb;
  wire [20:0] p3_add_33661_comb;
  wire [28:0] p3_add_33663_comb;
  wire [24:0] p3_add_33665_comb;
  wire [20:0] p3_add_33667_comb;
  wire [28:0] p3_add_33669_comb;
  wire [24:0] p3_add_33673_comb;
  wire [20:0] p3_add_33675_comb;
  wire [28:0] p3_add_33677_comb;
  wire [24:0] p3_add_33679_comb;
  wire [20:0] p3_add_33681_comb;
  wire [28:0] p3_add_33683_comb;
  wire [24:0] p3_add_33751_comb;
  wire [20:0] p3_add_33753_comb;
  wire [30:0] p3_add_33755_comb;
  wire [24:0] p3_add_33757_comb;
  wire [20:0] p3_add_33759_comb;
  wire [30:0] p3_add_33761_comb;
  wire [24:0] p3_add_33773_comb;
  wire [20:0] p3_add_33775_comb;
  wire [28:0] p3_add_33777_comb;
  wire [24:0] p3_add_33779_comb;
  wire [20:0] p3_add_33781_comb;
  wire [28:0] p3_add_33783_comb;
  wire [24:0] p3_add_33789_comb;
  wire [20:0] p3_add_33791_comb;
  wire [28:0] p3_add_33793_comb;
  wire [24:0] p3_add_33795_comb;
  wire [20:0] p3_add_33797_comb;
  wire [28:0] p3_add_33799_comb;
  wire [24:0] p3_add_33957_comb;
  wire [20:0] p3_add_33959_comb;
  wire [30:0] p3_add_33961_comb;
  wire [24:0] p3_add_33963_comb;
  wire [20:0] p3_add_33965_comb;
  wire [30:0] p3_add_33967_comb;
  wire [24:0] p3_add_33969_comb;
  wire [20:0] p3_add_33971_comb;
  wire [28:0] p3_add_33973_comb;
  wire [24:0] p3_add_33975_comb;
  wire [20:0] p3_add_33977_comb;
  wire [28:0] p3_add_33979_comb;
  wire [24:0] p3_add_33981_comb;
  wire [20:0] p3_add_33983_comb;
  wire [28:0] p3_add_33985_comb;
  wire [24:0] p3_add_33987_comb;
  wire [20:0] p3_add_33989_comb;
  wire [28:0] p3_add_33991_comb;
  wire [28:0] p3_add_33481_comb;
  wire [31:0] p3_add_33483_comb;
  wire [31:0] p3_add_33484_comb;
  wire [28:0] p3_add_33485_comb;
  wire [31:0] p3_add_33487_comb;
  wire [31:0] p3_add_33488_comb;
  wire [28:0] p3_add_33505_comb;
  wire [31:0] p3_add_33507_comb;
  wire [31:0] p3_add_33508_comb;
  wire [28:0] p3_add_33509_comb;
  wire [31:0] p3_add_33511_comb;
  wire [31:0] p3_add_33512_comb;
  wire [28:0] p3_add_33577_comb;
  wire [31:0] p3_add_33579_comb;
  wire [31:0] p3_add_33580_comb;
  wire [28:0] p3_add_33581_comb;
  wire [31:0] p3_add_33583_comb;
  wire [31:0] p3_add_33584_comb;
  wire [31:0] p3_sub_33689_comb;
  wire [31:0] p3_sub_33692_comb;
  wire [29:0] p3_concat_33710_comb;
  wire [29:0] p3_concat_33714_comb;
  wire [31:0] p3_sub_33807_comb;
  wire [31:0] p3_sub_33810_comb;
  wire [29:0] p3_concat_33820_comb;
  wire [29:0] p3_concat_33824_comb;
  wire [31:0] p3_sub_33993_comb;
  wire [31:0] p3_sub_33996_comb;
  wire [29:0] p3_concat_34002_comb;
  wire [29:0] p3_concat_34006_comb;
  wire [31:0] p3_add_33745_comb;
  wire [24:0] p3_add_33746_comb;
  wire [31:0] p3_add_33748_comb;
  wire [24:0] p3_add_33749_comb;
  wire [28:0] p3_add_33763_comb;
  wire [29:0] p3_add_33765_comb;
  wire [28:0] p3_add_33768_comb;
  wire [29:0] p3_add_33770_comb;
  wire [30:0] p3_add_33785_comb;
  wire [29:0] p3_add_33786_comb;
  wire [30:0] p3_add_33787_comb;
  wire [29:0] p3_add_33788_comb;
  wire [29:0] p3_add_33801_comb;
  wire [29:0] p3_add_33803_comb;
  wire [29:0] p3_add_33804_comb;
  wire [29:0] p3_add_33806_comb;
  wire [31:0] p3_add_33849_comb;
  wire [24:0] p3_add_33850_comb;
  wire [31:0] p3_add_33852_comb;
  wire [24:0] p3_add_33853_comb;
  wire [28:0] p3_add_33857_comb;
  wire [29:0] p3_add_33859_comb;
  wire [28:0] p3_add_33862_comb;
  wire [29:0] p3_add_33864_comb;
  wire [30:0] p3_add_33869_comb;
  wire [29:0] p3_add_33870_comb;
  wire [30:0] p3_add_33871_comb;
  wire [29:0] p3_add_33872_comb;
  wire [29:0] p3_add_33875_comb;
  wire [29:0] p3_add_33877_comb;
  wire [29:0] p3_add_33878_comb;
  wire [29:0] p3_add_33880_comb;
  wire [31:0] p3_add_34019_comb;
  wire [24:0] p3_add_34020_comb;
  wire [31:0] p3_add_34022_comb;
  wire [24:0] p3_add_34023_comb;
  wire [28:0] p3_add_34025_comb;
  wire [29:0] p3_add_34027_comb;
  wire [28:0] p3_add_34030_comb;
  wire [29:0] p3_add_34032_comb;
  wire [30:0] p3_add_34035_comb;
  wire [29:0] p3_add_34036_comb;
  wire [30:0] p3_add_34037_comb;
  wire [29:0] p3_add_34038_comb;
  wire [29:0] p3_add_34039_comb;
  wire [29:0] p3_add_34041_comb;
  wire [29:0] p3_add_34042_comb;
  wire [29:0] p3_add_34044_comb;
  wire [28:0] p3_add_33501_comb;
  wire [28:0] p3_add_33503_comb;
  wire [30:0] p3_add_33513_comb;
  wire [28:0] p3_add_33515_comb;
  wire [30:0] p3_add_33517_comb;
  wire [28:0] p3_add_33519_comb;
  wire [28:0] p3_add_33535_comb;
  wire [28:0] p3_add_33537_comb;
  wire [30:0] p3_add_33541_comb;
  wire [28:0] p3_add_33543_comb;
  wire [30:0] p3_add_33545_comb;
  wire [28:0] p3_add_33547_comb;
  wire [28:0] p3_add_33595_comb;
  wire [28:0] p3_add_33597_comb;
  wire [30:0] p3_add_33599_comb;
  wire [28:0] p3_add_33601_comb;
  wire [30:0] p3_add_33603_comb;
  wire [28:0] p3_add_33605_comb;
  wire [31:0] p3_add_33521_comb;
  wire [31:0] p3_add_33523_comb;
  wire [31:0] p3_add_33555_comb;
  wire [31:0] p3_add_33557_comb;
  wire [31:0] p3_add_33637_comb;
  wire [31:0] p3_add_33639_comb;
  wire [29:0] p3_add_33855_comb;
  wire [29:0] p3_add_33856_comb;
  wire [31:0] p3_sub_33867_comb;
  wire [31:0] p3_sub_33868_comb;
  wire [31:0] p3_sub_33873_comb;
  wire [31:0] p3_sub_33874_comb;
  wire [31:0] p3_sub_33881_comb;
  wire [31:0] p3_sub_33882_comb;
  wire [29:0] p3_add_33911_comb;
  wire [29:0] p3_add_33912_comb;
  wire [31:0] p3_sub_33913_comb;
  wire [31:0] p3_sub_33914_comb;
  wire [31:0] p3_sub_33915_comb;
  wire [31:0] p3_sub_33916_comb;
  wire [31:0] p3_sub_33917_comb;
  wire [31:0] p3_sub_33918_comb;
  wire [29:0] p3_add_34061_comb;
  wire [29:0] p3_add_34062_comb;
  wire [31:0] p3_sub_34063_comb;
  wire [31:0] p3_sub_34064_comb;
  wire [31:0] p3_sub_34065_comb;
  wire [31:0] p3_sub_34066_comb;
  wire [31:0] p3_sub_34067_comb;
  wire [31:0] p3_sub_34068_comb;
  wire [31:0] p3_sub_33539_comb;
  wire [31:0] p3_sub_33540_comb;
  wire [31:0] p3_sub_33549_comb;
  wire [31:0] p3_sub_33550_comb;
  wire [31:0] p3_sub_33567_comb;
  wire [31:0] p3_sub_33568_comb;
  wire [31:0] p3_sub_33569_comb;
  wire [31:0] p3_sub_33570_comb;
  wire [31:0] p3_sub_33685_comb;
  wire [31:0] p3_sub_33686_comb;
  wire [31:0] p3_sub_33687_comb;
  wire [31:0] p3_sub_33688_comb;
  wire [23:0] p3_bit_slice_33889_comb;
  wire [23:0] p3_bit_slice_33890_comb;
  wire [23:0] p3_bit_slice_33895_comb;
  wire [23:0] p3_bit_slice_33896_comb;
  wire [23:0] p3_bit_slice_33901_comb;
  wire [23:0] p3_bit_slice_33902_comb;
  wire [23:0] p3_bit_slice_33907_comb;
  wire [23:0] p3_bit_slice_33908_comb;
  wire [23:0] p3_bit_slice_33947_comb;
  wire [23:0] p3_bit_slice_33948_comb;
  wire [23:0] p3_bit_slice_33949_comb;
  wire [23:0] p3_bit_slice_33950_comb;
  wire [23:0] p3_bit_slice_33951_comb;
  wire [23:0] p3_bit_slice_33952_comb;
  wire [23:0] p3_bit_slice_33953_comb;
  wire [23:0] p3_bit_slice_33954_comb;
  wire [23:0] p3_bit_slice_34069_comb;
  wire [23:0] p3_bit_slice_34070_comb;
  wire [23:0] p3_bit_slice_34071_comb;
  wire [23:0] p3_bit_slice_34072_comb;
  wire [23:0] p3_bit_slice_34073_comb;
  wire [23:0] p3_bit_slice_34074_comb;
  wire [23:0] p3_bit_slice_34075_comb;
  wire [23:0] p3_bit_slice_34076_comb;
  assign p3_add_33593_comb = p2_bit_slice_33265 + p2_umul_33254[31:5];
  assign p3_add_33594_comb = p2_bit_slice_33266 + p2_umul_33256[31:5];
  assign p3_add_33671_comb = p2_bit_slice_33275 + p2_umul_33270[31:5];
  assign p3_add_33672_comb = p2_bit_slice_33276 + p2_umul_33272[31:5];
  assign p3_add_33909_comb = p2_bit_slice_33291 + p2_umul_33286[31:5];
  assign p3_add_33910_comb = p2_bit_slice_33292 + p2_umul_33288[31:5];
  assign p3_add_33463_comb = p2_umul_33169[31:2] + p2_umul_33170[31:2];
  assign p3_add_33465_comb = p2_umul_33171[31:2] + p2_umul_33172[31:2];
  assign p3_add_33477_comb = p2_umul_33185[31:2] + p2_umul_33186[31:2];
  assign p3_add_33479_comb = p2_umul_33187[31:2] + p2_umul_33188[31:2];
  assign p3_add_33563_comb = p2_umul_33225[31:2] + p2_umul_33226[31:2];
  assign p3_add_33565_comb = p2_umul_33227[31:2] + p2_umul_33228[31:2];
  assign p3_add_33610_comb = p2_bit_slice_32973 + p2_bit_slice_32974;
  assign p3_add_33616_comb = p2_bit_slice_32975 + p2_bit_slice_32976;
  assign p3_add_33698_comb = p2_bit_slice_32989 + p2_bit_slice_32990;
  assign p3_add_33704_comb = p2_bit_slice_32991 + p2_bit_slice_32992;
  assign p3_add_33922_comb = p2_bit_slice_33011 + p2_bit_slice_33012;
  assign p3_add_33928_comb = p2_bit_slice_33013 + p2_bit_slice_33014;
  assign p3_concat_33473_comb = {p3_add_33463_comb, p2_umul_33170[1:0]};
  assign p3_concat_33476_comb = {p3_add_33465_comb, p2_umul_33172[1:0]};
  assign p3_concat_33491_comb = {p3_add_33477_comb, p2_umul_33186[1:0]};
  assign p3_concat_33494_comb = {p3_add_33479_comb, p2_umul_33188[1:0]};
  assign p3_concat_33573_comb = {p3_add_33563_comb, p2_umul_33226[1:0]};
  assign p3_concat_33576_comb = {p3_add_33565_comb, p2_umul_33228[1:0]};
  assign p3_add_33647_comb = p2_umul_33189[31:7] + 25'h000_0001;
  assign p3_add_33649_comb = p2_umul_33170[31:11] + p3_add_33610_comb;
  assign p3_add_33651_comb = p2_umul_33204[31:1] + p2_umul_33190[31:1];
  assign p3_add_33653_comb = p2_umul_33193[31:7] + 25'h000_0001;
  assign p3_add_33655_comb = p2_umul_33172[31:11] + p3_add_33616_comb;
  assign p3_add_33657_comb = p2_umul_33206[31:1] + p2_umul_33194[31:1];
  assign p3_add_33659_comb = p2_umul_33204[31:7] + 25'h000_0001;
  assign p3_add_33661_comb = p2_umul_33190[31:11] + p3_add_33610_comb;
  assign p3_add_33663_comb = p2_umul_33189[31:3] + p2_umul_33170[31:3];
  assign p3_add_33665_comb = p2_umul_33206[31:7] + 25'h000_0001;
  assign p3_add_33667_comb = p2_umul_33194[31:11] + p3_add_33616_comb;
  assign p3_add_33669_comb = p2_umul_33193[31:3] + p2_umul_33172[31:3];
  assign p3_add_33673_comb = p2_umul_33203[31:7] + 25'h000_0001;
  assign p3_add_33675_comb = p3_add_33593_comb[26:6] + p3_add_33610_comb;
  assign p3_add_33677_comb = p2_umul_33189[31:3] + p2_umul_33169[31:3];
  assign p3_add_33679_comb = p2_umul_33205[31:7] + 25'h000_0001;
  assign p3_add_33681_comb = p3_add_33594_comb[26:6] + p3_add_33616_comb;
  assign p3_add_33683_comb = p2_umul_33193[31:3] + p2_umul_33171[31:3];
  assign p3_add_33751_comb = p2_umul_33207[31:7] + 25'h000_0001;
  assign p3_add_33753_comb = p2_umul_33186[31:11] + p3_add_33698_comb;
  assign p3_add_33755_comb = p2_umul_33216[31:1] + p2_umul_33208[31:1];
  assign p3_add_33757_comb = p2_umul_33211[31:7] + 25'h000_0001;
  assign p3_add_33759_comb = p2_umul_33188[31:11] + p3_add_33704_comb;
  assign p3_add_33761_comb = p2_umul_33218[31:1] + p2_umul_33212[31:1];
  assign p3_add_33773_comb = p2_umul_33216[31:7] + 25'h000_0001;
  assign p3_add_33775_comb = p2_umul_33208[31:11] + p3_add_33698_comb;
  assign p3_add_33777_comb = p2_umul_33207[31:3] + p2_umul_33186[31:3];
  assign p3_add_33779_comb = p2_umul_33218[31:7] + 25'h000_0001;
  assign p3_add_33781_comb = p2_umul_33212[31:11] + p3_add_33704_comb;
  assign p3_add_33783_comb = p2_umul_33211[31:3] + p2_umul_33188[31:3];
  assign p3_add_33789_comb = p2_umul_33215[31:7] + 25'h000_0001;
  assign p3_add_33791_comb = p3_add_33671_comb[26:6] + p3_add_33698_comb;
  assign p3_add_33793_comb = p2_umul_33207[31:3] + p2_umul_33185[31:3];
  assign p3_add_33795_comb = p2_umul_33217[31:7] + 25'h000_0001;
  assign p3_add_33797_comb = p3_add_33672_comb[26:6] + p3_add_33704_comb;
  assign p3_add_33799_comb = p2_umul_33211[31:3] + p2_umul_33187[31:3];
  assign p3_add_33957_comb = p2_umul_33235[31:7] + 25'h000_0001;
  assign p3_add_33959_comb = p2_umul_33226[31:11] + p3_add_33922_comb;
  assign p3_add_33961_comb = p2_umul_33250[31:1] + p2_umul_33236[31:1];
  assign p3_add_33963_comb = p2_umul_33239[31:7] + 25'h000_0001;
  assign p3_add_33965_comb = p2_umul_33228[31:11] + p3_add_33928_comb;
  assign p3_add_33967_comb = p2_umul_33252[31:1] + p2_umul_33240[31:1];
  assign p3_add_33969_comb = p2_umul_33250[31:7] + 25'h000_0001;
  assign p3_add_33971_comb = p2_umul_33236[31:11] + p3_add_33922_comb;
  assign p3_add_33973_comb = p2_umul_33235[31:3] + p2_umul_33226[31:3];
  assign p3_add_33975_comb = p2_umul_33252[31:7] + 25'h000_0001;
  assign p3_add_33977_comb = p2_umul_33240[31:11] + p3_add_33928_comb;
  assign p3_add_33979_comb = p2_umul_33239[31:3] + p2_umul_33228[31:3];
  assign p3_add_33981_comb = p2_umul_33249[31:7] + 25'h000_0001;
  assign p3_add_33983_comb = p3_add_33909_comb[26:6] + p3_add_33922_comb;
  assign p3_add_33985_comb = p2_umul_33235[31:3] + p2_umul_33225[31:3];
  assign p3_add_33987_comb = p2_umul_33251[31:7] + 25'h000_0001;
  assign p3_add_33989_comb = p3_add_33910_comb[26:6] + p3_add_33928_comb;
  assign p3_add_33991_comb = p2_umul_33239[31:3] + p2_umul_33227[31:3];
  assign p3_add_33481_comb = p2_umul_33189[31:3] + p2_umul_33190[31:3];
  assign p3_add_33483_comb = p2_umul_33203 + p3_concat_33473_comb;
  assign p3_add_33484_comb = p2_umul_33204 + p2_umul_33170;
  assign p3_add_33485_comb = p2_umul_33193[31:3] + p2_umul_33194[31:3];
  assign p3_add_33487_comb = p2_umul_33205 + p3_concat_33476_comb;
  assign p3_add_33488_comb = p2_umul_33206 + p2_umul_33172;
  assign p3_add_33505_comb = p2_umul_33207[31:3] + p2_umul_33208[31:3];
  assign p3_add_33507_comb = p2_umul_33215 + p3_concat_33491_comb;
  assign p3_add_33508_comb = p2_umul_33216 + p2_umul_33186;
  assign p3_add_33509_comb = p2_umul_33211[31:3] + p2_umul_33212[31:3];
  assign p3_add_33511_comb = p2_umul_33217 + p3_concat_33494_comb;
  assign p3_add_33512_comb = p2_umul_33218 + p2_umul_33188;
  assign p3_add_33577_comb = p2_umul_33235[31:3] + p2_umul_33236[31:3];
  assign p3_add_33579_comb = p2_umul_33249 + p3_concat_33573_comb;
  assign p3_add_33580_comb = p2_umul_33250 + p2_umul_33226;
  assign p3_add_33581_comb = p2_umul_33239[31:3] + p2_umul_33240[31:3];
  assign p3_add_33583_comb = p2_umul_33251 + p3_concat_33576_comb;
  assign p3_add_33584_comb = p2_umul_33252 + p2_umul_33228;
  assign p3_sub_33689_comb = p2_umul_33189 - p2_umul_33203;
  assign p3_sub_33692_comb = p2_umul_33193 - p2_umul_33205;
  assign p3_concat_33710_comb = {p3_add_33593_comb, p2_umul_33254[4:2]};
  assign p3_concat_33714_comb = {p3_add_33594_comb, p2_umul_33256[4:2]};
  assign p3_sub_33807_comb = p2_umul_33207 - p2_umul_33215;
  assign p3_sub_33810_comb = p2_umul_33211 - p2_umul_33217;
  assign p3_concat_33820_comb = {p3_add_33671_comb, p2_umul_33270[4:2]};
  assign p3_concat_33824_comb = {p3_add_33672_comb, p2_umul_33272[4:2]};
  assign p3_sub_33993_comb = p2_umul_33235 - p2_umul_33249;
  assign p3_sub_33996_comb = p2_umul_33239 - p2_umul_33251;
  assign p3_concat_34002_comb = {p3_add_33909_comb, p2_umul_33286[4:2]};
  assign p3_concat_34006_comb = {p3_add_33910_comb, p2_umul_33288[4:2]};
  assign p3_add_33745_comb = p3_sub_33689_comb + p3_concat_33473_comb;
  assign p3_add_33746_comb = p3_add_33593_comb[26:2] + {p3_add_33610_comb, 4'h1};
  assign p3_add_33748_comb = p3_sub_33692_comb + p3_concat_33476_comb;
  assign p3_add_33749_comb = p3_add_33594_comb[26:2] + {p3_add_33616_comb, 4'h1};
  assign p3_add_33763_comb = {p3_add_33647_comb, p2_umul_33189[6:3]} + {p3_add_33649_comb, p2_umul_33170[10:3]};
  assign p3_add_33765_comb = p3_add_33651_comb[30:1] + p3_concat_33710_comb;
  assign p3_add_33768_comb = {p3_add_33653_comb, p2_umul_33193[6:3]} + {p3_add_33655_comb, p2_umul_33172[10:3]};
  assign p3_add_33770_comb = p3_add_33657_comb[30:1] + p3_concat_33714_comb;
  assign p3_add_33785_comb = {p3_add_33659_comb, p2_umul_33204[6:1]} + {p3_add_33661_comb, p2_umul_33190[10:1]};
  assign p3_add_33786_comb = {p3_add_33663_comb, p2_umul_33170[2]} + p3_concat_33710_comb;
  assign p3_add_33787_comb = {p3_add_33665_comb, p2_umul_33206[6:1]} + {p3_add_33667_comb, p2_umul_33194[10:1]};
  assign p3_add_33788_comb = {p3_add_33669_comb, p2_umul_33172[2]} + p3_concat_33714_comb;
  assign p3_add_33801_comb = {p3_add_33673_comb, p2_umul_33203[6:2]} + {p3_add_33675_comb, p3_add_33593_comb[5:0], p2_umul_33254[4:2]};
  assign p3_add_33803_comb = {p3_add_33677_comb, p2_umul_33169[2]} + p2_umul_33170[31:2];
  assign p3_add_33804_comb = {p3_add_33679_comb, p2_umul_33205[6:2]} + {p3_add_33681_comb, p3_add_33594_comb[5:0], p2_umul_33256[4:2]};
  assign p3_add_33806_comb = {p3_add_33683_comb, p2_umul_33171[2]} + p2_umul_33172[31:2];
  assign p3_add_33849_comb = p3_sub_33807_comb + p3_concat_33491_comb;
  assign p3_add_33850_comb = p3_add_33671_comb[26:2] + {p3_add_33698_comb, 4'h1};
  assign p3_add_33852_comb = p3_sub_33810_comb + p3_concat_33494_comb;
  assign p3_add_33853_comb = p3_add_33672_comb[26:2] + {p3_add_33704_comb, 4'h1};
  assign p3_add_33857_comb = {p3_add_33751_comb, p2_umul_33207[6:3]} + {p3_add_33753_comb, p2_umul_33186[10:3]};
  assign p3_add_33859_comb = p3_add_33755_comb[30:1] + p3_concat_33820_comb;
  assign p3_add_33862_comb = {p3_add_33757_comb, p2_umul_33211[6:3]} + {p3_add_33759_comb, p2_umul_33188[10:3]};
  assign p3_add_33864_comb = p3_add_33761_comb[30:1] + p3_concat_33824_comb;
  assign p3_add_33869_comb = {p3_add_33773_comb, p2_umul_33216[6:1]} + {p3_add_33775_comb, p2_umul_33208[10:1]};
  assign p3_add_33870_comb = {p3_add_33777_comb, p2_umul_33186[2]} + p3_concat_33820_comb;
  assign p3_add_33871_comb = {p3_add_33779_comb, p2_umul_33218[6:1]} + {p3_add_33781_comb, p2_umul_33212[10:1]};
  assign p3_add_33872_comb = {p3_add_33783_comb, p2_umul_33188[2]} + p3_concat_33824_comb;
  assign p3_add_33875_comb = {p3_add_33789_comb, p2_umul_33215[6:2]} + {p3_add_33791_comb, p3_add_33671_comb[5:0], p2_umul_33270[4:2]};
  assign p3_add_33877_comb = {p3_add_33793_comb, p2_umul_33185[2]} + p2_umul_33186[31:2];
  assign p3_add_33878_comb = {p3_add_33795_comb, p2_umul_33217[6:2]} + {p3_add_33797_comb, p3_add_33672_comb[5:0], p2_umul_33272[4:2]};
  assign p3_add_33880_comb = {p3_add_33799_comb, p2_umul_33187[2]} + p2_umul_33188[31:2];
  assign p3_add_34019_comb = p3_sub_33993_comb + p3_concat_33573_comb;
  assign p3_add_34020_comb = p3_add_33909_comb[26:2] + {p3_add_33922_comb, 4'h1};
  assign p3_add_34022_comb = p3_sub_33996_comb + p3_concat_33576_comb;
  assign p3_add_34023_comb = p3_add_33910_comb[26:2] + {p3_add_33928_comb, 4'h1};
  assign p3_add_34025_comb = {p3_add_33957_comb, p2_umul_33235[6:3]} + {p3_add_33959_comb, p2_umul_33226[10:3]};
  assign p3_add_34027_comb = p3_add_33961_comb[30:1] + p3_concat_34002_comb;
  assign p3_add_34030_comb = {p3_add_33963_comb, p2_umul_33239[6:3]} + {p3_add_33965_comb, p2_umul_33228[10:3]};
  assign p3_add_34032_comb = p3_add_33967_comb[30:1] + p3_concat_34006_comb;
  assign p3_add_34035_comb = {p3_add_33969_comb, p2_umul_33250[6:1]} + {p3_add_33971_comb, p2_umul_33236[10:1]};
  assign p3_add_34036_comb = {p3_add_33973_comb, p2_umul_33226[2]} + p3_concat_34002_comb;
  assign p3_add_34037_comb = {p3_add_33975_comb, p2_umul_33252[6:1]} + {p3_add_33977_comb, p2_umul_33240[10:1]};
  assign p3_add_34038_comb = {p3_add_33979_comb, p2_umul_33228[2]} + p3_concat_34006_comb;
  assign p3_add_34039_comb = {p3_add_33981_comb, p2_umul_33249[6:2]} + {p3_add_33983_comb, p3_add_33909_comb[5:0], p2_umul_33286[4:2]};
  assign p3_add_34041_comb = {p3_add_33985_comb, p2_umul_33225[2]} + p2_umul_33226[31:2];
  assign p3_add_34042_comb = {p3_add_33987_comb, p2_umul_33251[6:2]} + {p3_add_33989_comb, p3_add_33910_comb[5:0], p2_umul_33288[4:2]};
  assign p3_add_34044_comb = {p3_add_33991_comb, p2_umul_33227[2]} + p2_umul_33228[31:2];
  assign p3_add_33501_comb = p3_add_33481_comb + p2_umul_33189[31:3];
  assign p3_add_33503_comb = p3_add_33485_comb + p2_umul_33193[31:3];
  assign p3_add_33513_comb = {p3_add_33481_comb, p2_umul_33190[2:1]} + p3_add_33483_comb[31:1];
  assign p3_add_33515_comb = p3_add_33484_comb[31:3] + p2_umul_33189[31:3];
  assign p3_add_33517_comb = {p3_add_33485_comb, p2_umul_33194[2:1]} + p3_add_33487_comb[31:1];
  assign p3_add_33519_comb = p3_add_33488_comb[31:3] + p2_umul_33193[31:3];
  assign p3_add_33535_comb = p3_add_33505_comb + p2_umul_33207[31:3];
  assign p3_add_33537_comb = p3_add_33509_comb + p2_umul_33211[31:3];
  assign p3_add_33541_comb = {p3_add_33505_comb, p2_umul_33208[2:1]} + p3_add_33507_comb[31:1];
  assign p3_add_33543_comb = p3_add_33508_comb[31:3] + p2_umul_33207[31:3];
  assign p3_add_33545_comb = {p3_add_33509_comb, p2_umul_33212[2:1]} + p3_add_33511_comb[31:1];
  assign p3_add_33547_comb = p3_add_33512_comb[31:3] + p2_umul_33211[31:3];
  assign p3_add_33595_comb = p3_add_33577_comb + p2_umul_33235[31:3];
  assign p3_add_33597_comb = p3_add_33581_comb + p2_umul_33239[31:3];
  assign p3_add_33599_comb = {p3_add_33577_comb, p2_umul_33236[2:1]} + p3_add_33579_comb[31:1];
  assign p3_add_33601_comb = p3_add_33580_comb[31:3] + p2_umul_33235[31:3];
  assign p3_add_33603_comb = {p3_add_33581_comb, p2_umul_33240[2:1]} + p3_add_33583_comb[31:1];
  assign p3_add_33605_comb = p3_add_33584_comb[31:3] + p2_umul_33239[31:3];
  assign p3_add_33521_comb = p3_add_33483_comb + p3_add_33484_comb;
  assign p3_add_33523_comb = p3_add_33487_comb + p3_add_33488_comb;
  assign p3_add_33555_comb = p3_add_33507_comb + p3_add_33508_comb;
  assign p3_add_33557_comb = p3_add_33511_comb + p3_add_33512_comb;
  assign p3_add_33637_comb = p3_add_33579_comb + p3_add_33580_comb;
  assign p3_add_33639_comb = p3_add_33583_comb + p3_add_33584_comb;
  assign p3_add_33855_comb = p3_add_33745_comb[31:2] + {p3_add_33746_comb, p3_add_33593_comb[1:0], p2_umul_33254[4:2]};
  assign p3_add_33856_comb = p3_add_33748_comb[31:2] + {p3_add_33749_comb, p3_add_33594_comb[1:0], p2_umul_33256[4:2]};
  assign p3_sub_33867_comb = {p3_add_33763_comb, p2_umul_33170[2:0]} - {p3_add_33765_comb, p3_add_33651_comb[0], p2_umul_33204[0]};
  assign p3_sub_33868_comb = {p3_add_33768_comb, p2_umul_33172[2:0]} - {p3_add_33770_comb, p3_add_33657_comb[0], p2_umul_33206[0]};
  assign p3_sub_33873_comb = {p3_add_33785_comb, p2_umul_33204[0]} - {p3_add_33786_comb, p2_umul_33170[1:0]};
  assign p3_sub_33874_comb = {p3_add_33787_comb, p2_umul_33206[0]} - {p3_add_33788_comb, p2_umul_33172[1:0]};
  assign p3_sub_33881_comb = {p3_add_33801_comb, p2_umul_33203[1:0]} - {p3_add_33803_comb, p2_umul_33170[1:0]};
  assign p3_sub_33882_comb = {p3_add_33804_comb, p2_umul_33205[1:0]} - {p3_add_33806_comb, p2_umul_33172[1:0]};
  assign p3_add_33911_comb = p3_add_33849_comb[31:2] + {p3_add_33850_comb, p3_add_33671_comb[1:0], p2_umul_33270[4:2]};
  assign p3_add_33912_comb = p3_add_33852_comb[31:2] + {p3_add_33853_comb, p3_add_33672_comb[1:0], p2_umul_33272[4:2]};
  assign p3_sub_33913_comb = {p3_add_33857_comb, p2_umul_33186[2:0]} - {p3_add_33859_comb, p3_add_33755_comb[0], p2_umul_33216[0]};
  assign p3_sub_33914_comb = {p3_add_33862_comb, p2_umul_33188[2:0]} - {p3_add_33864_comb, p3_add_33761_comb[0], p2_umul_33218[0]};
  assign p3_sub_33915_comb = {p3_add_33869_comb, p2_umul_33216[0]} - {p3_add_33870_comb, p2_umul_33186[1:0]};
  assign p3_sub_33916_comb = {p3_add_33871_comb, p2_umul_33218[0]} - {p3_add_33872_comb, p2_umul_33188[1:0]};
  assign p3_sub_33917_comb = {p3_add_33875_comb, p2_umul_33215[1:0]} - {p3_add_33877_comb, p2_umul_33186[1:0]};
  assign p3_sub_33918_comb = {p3_add_33878_comb, p2_umul_33217[1:0]} - {p3_add_33880_comb, p2_umul_33188[1:0]};
  assign p3_add_34061_comb = p3_add_34019_comb[31:2] + {p3_add_34020_comb, p3_add_33909_comb[1:0], p2_umul_33286[4:2]};
  assign p3_add_34062_comb = p3_add_34022_comb[31:2] + {p3_add_34023_comb, p3_add_33910_comb[1:0], p2_umul_33288[4:2]};
  assign p3_sub_34063_comb = {p3_add_34025_comb, p2_umul_33226[2:0]} - {p3_add_34027_comb, p3_add_33961_comb[0], p2_umul_33250[0]};
  assign p3_sub_34064_comb = {p3_add_34030_comb, p2_umul_33228[2:0]} - {p3_add_34032_comb, p3_add_33967_comb[0], p2_umul_33252[0]};
  assign p3_sub_34065_comb = {p3_add_34035_comb, p2_umul_33250[0]} - {p3_add_34036_comb, p2_umul_33226[1:0]};
  assign p3_sub_34066_comb = {p3_add_34037_comb, p2_umul_33252[0]} - {p3_add_34038_comb, p2_umul_33228[1:0]};
  assign p3_sub_34067_comb = {p3_add_34039_comb, p2_umul_33249[1:0]} - {p3_add_34041_comb, p2_umul_33226[1:0]};
  assign p3_sub_34068_comb = {p3_add_34042_comb, p2_umul_33251[1:0]} - {p3_add_34044_comb, p2_umul_33228[1:0]};
  assign p3_sub_33539_comb = p3_add_33521_comb - {p3_add_33501_comb, p2_umul_33190[2:0]};
  assign p3_sub_33540_comb = p3_add_33523_comb - {p3_add_33503_comb, p2_umul_33194[2:0]};
  assign p3_sub_33549_comb = {p3_add_33513_comb, p3_add_33483_comb[0]} - {p3_add_33515_comb, p3_add_33484_comb[2:0]};
  assign p3_sub_33550_comb = {p3_add_33517_comb, p3_add_33487_comb[0]} - {p3_add_33519_comb, p3_add_33488_comb[2:0]};
  assign p3_sub_33567_comb = p3_add_33555_comb - {p3_add_33535_comb, p2_umul_33208[2:0]};
  assign p3_sub_33568_comb = p3_add_33557_comb - {p3_add_33537_comb, p2_umul_33212[2:0]};
  assign p3_sub_33569_comb = {p3_add_33541_comb, p3_add_33507_comb[0]} - {p3_add_33543_comb, p3_add_33508_comb[2:0]};
  assign p3_sub_33570_comb = {p3_add_33545_comb, p3_add_33511_comb[0]} - {p3_add_33547_comb, p3_add_33512_comb[2:0]};
  assign p3_sub_33685_comb = p3_add_33637_comb - {p3_add_33595_comb, p2_umul_33236[2:0]};
  assign p3_sub_33686_comb = p3_add_33639_comb - {p3_add_33597_comb, p2_umul_33240[2:0]};
  assign p3_sub_33687_comb = {p3_add_33599_comb, p3_add_33579_comb[0]} - {p3_add_33601_comb, p3_add_33580_comb[2:0]};
  assign p3_sub_33688_comb = {p3_add_33603_comb, p3_add_33583_comb[0]} - {p3_add_33605_comb, p3_add_33584_comb[2:0]};
  assign p3_bit_slice_33889_comb = p3_add_33855_comb[29:6];
  assign p3_bit_slice_33890_comb = p3_add_33856_comb[29:6];
  assign p3_bit_slice_33895_comb = p3_sub_33867_comb[31:8];
  assign p3_bit_slice_33896_comb = p3_sub_33868_comb[31:8];
  assign p3_bit_slice_33901_comb = p3_sub_33873_comb[31:8];
  assign p3_bit_slice_33902_comb = p3_sub_33874_comb[31:8];
  assign p3_bit_slice_33907_comb = p3_sub_33881_comb[31:8];
  assign p3_bit_slice_33908_comb = p3_sub_33882_comb[31:8];
  assign p3_bit_slice_33947_comb = p3_add_33911_comb[29:6];
  assign p3_bit_slice_33948_comb = p3_add_33912_comb[29:6];
  assign p3_bit_slice_33949_comb = p3_sub_33913_comb[31:8];
  assign p3_bit_slice_33950_comb = p3_sub_33914_comb[31:8];
  assign p3_bit_slice_33951_comb = p3_sub_33915_comb[31:8];
  assign p3_bit_slice_33952_comb = p3_sub_33916_comb[31:8];
  assign p3_bit_slice_33953_comb = p3_sub_33917_comb[31:8];
  assign p3_bit_slice_33954_comb = p3_sub_33918_comb[31:8];
  assign p3_bit_slice_34069_comb = p3_add_34061_comb[29:6];
  assign p3_bit_slice_34070_comb = p3_add_34062_comb[29:6];
  assign p3_bit_slice_34071_comb = p3_sub_34063_comb[31:8];
  assign p3_bit_slice_34072_comb = p3_sub_34064_comb[31:8];
  assign p3_bit_slice_34073_comb = p3_sub_34065_comb[31:8];
  assign p3_bit_slice_34074_comb = p3_sub_34066_comb[31:8];
  assign p3_bit_slice_34075_comb = p3_sub_34067_comb[31:8];
  assign p3_bit_slice_34076_comb = p3_sub_34068_comb[31:8];

  // Registers for pipe stage 3:
  reg [31:0] p3_sub_33539;
  reg [31:0] p3_sub_33540;
  reg [31:0] p3_sub_33549;
  reg [31:0] p3_sub_33550;
  reg [31:0] p3_sub_33567;
  reg [31:0] p3_sub_33568;
  reg [31:0] p3_sub_33569;
  reg [31:0] p3_sub_33570;
  reg [31:0] p3_array_index_32965;
  reg [31:0] p3_array_index_32966;
  reg [20:0] p3_bit_slice_32973;
  reg [20:0] p3_bit_slice_32974;
  reg [20:0] p3_bit_slice_32975;
  reg [20:0] p3_bit_slice_32976;
  reg [31:0] p3_array_index_32979;
  reg [31:0] p3_array_index_32980;
  reg [31:0] p3_array_index_32985;
  reg [31:0] p3_array_index_32986;
  reg [20:0] p3_bit_slice_32989;
  reg [20:0] p3_bit_slice_32990;
  reg [20:0] p3_bit_slice_32991;
  reg [20:0] p3_bit_slice_32992;
  reg [31:0] p3_sub_33685;
  reg [31:0] p3_sub_33686;
  reg [31:0] p3_sub_33687;
  reg [31:0] p3_sub_33688;
  reg [31:0] p3_array_index_32997;
  reg [31:0] p3_array_index_32998;
  reg [23:0] p3_bit_slice_33889;
  reg [23:0] p3_bit_slice_33890;
  reg [23:0] p3_bit_slice_33895;
  reg [23:0] p3_bit_slice_33896;
  reg [23:0] p3_bit_slice_33901;
  reg [23:0] p3_bit_slice_33902;
  reg [23:0] p3_bit_slice_33907;
  reg [23:0] p3_bit_slice_33908;
  reg [20:0] p3_bit_slice_33011;
  reg [20:0] p3_bit_slice_33012;
  reg [20:0] p3_bit_slice_33013;
  reg [20:0] p3_bit_slice_33014;
  reg [23:0] p3_bit_slice_33947;
  reg [23:0] p3_bit_slice_33948;
  reg [23:0] p3_bit_slice_33949;
  reg [23:0] p3_bit_slice_33950;
  reg [23:0] p3_bit_slice_33951;
  reg [23:0] p3_bit_slice_33952;
  reg [23:0] p3_bit_slice_33953;
  reg [23:0] p3_bit_slice_33954;
  reg [31:0] p3_array_index_33017;
  reg [31:0] p3_array_index_33018;
  reg [31:0] p3_array_index_33021;
  reg [31:0] p3_array_index_33022;
  reg [23:0] p3_bit_slice_34069;
  reg [23:0] p3_bit_slice_34070;
  reg [23:0] p3_bit_slice_34071;
  reg [23:0] p3_bit_slice_34072;
  reg [23:0] p3_bit_slice_34073;
  reg [23:0] p3_bit_slice_34074;
  reg [23:0] p3_bit_slice_34075;
  reg [23:0] p3_bit_slice_34076;
  reg [20:0] p3_bit_slice_33029;
  reg [20:0] p3_bit_slice_33030;
  reg [20:0] p3_bit_slice_33033;
  reg [20:0] p3_bit_slice_33034;
  reg [31:0] p3_umul_33254;
  reg [31:0] p3_umul_33256;
  reg [31:0] p3_umul_33267;
  reg [31:0] p3_umul_33268;
  reg [31:0] p3_umul_33270;
  reg [31:0] p3_umul_33272;
  reg [31:0] p3_umul_33277;
  reg [31:0] p3_umul_33278;
  reg [31:0] p3_umul_33286;
  reg [31:0] p3_umul_33288;
  reg [31:0] p3_umul_33293;
  reg [31:0] p3_umul_33294;
  always_ff @ (posedge clk) begin
    p3_sub_33539 <= p3_sub_33539_comb;
    p3_sub_33540 <= p3_sub_33540_comb;
    p3_sub_33549 <= p3_sub_33549_comb;
    p3_sub_33550 <= p3_sub_33550_comb;
    p3_sub_33567 <= p3_sub_33567_comb;
    p3_sub_33568 <= p3_sub_33568_comb;
    p3_sub_33569 <= p3_sub_33569_comb;
    p3_sub_33570 <= p3_sub_33570_comb;
    p3_array_index_32965 <= p2_array_index_32965;
    p3_array_index_32966 <= p2_array_index_32966;
    p3_bit_slice_32973 <= p2_bit_slice_32973;
    p3_bit_slice_32974 <= p2_bit_slice_32974;
    p3_bit_slice_32975 <= p2_bit_slice_32975;
    p3_bit_slice_32976 <= p2_bit_slice_32976;
    p3_array_index_32979 <= p2_array_index_32979;
    p3_array_index_32980 <= p2_array_index_32980;
    p3_array_index_32985 <= p2_array_index_32985;
    p3_array_index_32986 <= p2_array_index_32986;
    p3_bit_slice_32989 <= p2_bit_slice_32989;
    p3_bit_slice_32990 <= p2_bit_slice_32990;
    p3_bit_slice_32991 <= p2_bit_slice_32991;
    p3_bit_slice_32992 <= p2_bit_slice_32992;
    p3_sub_33685 <= p3_sub_33685_comb;
    p3_sub_33686 <= p3_sub_33686_comb;
    p3_sub_33687 <= p3_sub_33687_comb;
    p3_sub_33688 <= p3_sub_33688_comb;
    p3_array_index_32997 <= p2_array_index_32997;
    p3_array_index_32998 <= p2_array_index_32998;
    p3_bit_slice_33889 <= p3_bit_slice_33889_comb;
    p3_bit_slice_33890 <= p3_bit_slice_33890_comb;
    p3_bit_slice_33895 <= p3_bit_slice_33895_comb;
    p3_bit_slice_33896 <= p3_bit_slice_33896_comb;
    p3_bit_slice_33901 <= p3_bit_slice_33901_comb;
    p3_bit_slice_33902 <= p3_bit_slice_33902_comb;
    p3_bit_slice_33907 <= p3_bit_slice_33907_comb;
    p3_bit_slice_33908 <= p3_bit_slice_33908_comb;
    p3_bit_slice_33011 <= p2_bit_slice_33011;
    p3_bit_slice_33012 <= p2_bit_slice_33012;
    p3_bit_slice_33013 <= p2_bit_slice_33013;
    p3_bit_slice_33014 <= p2_bit_slice_33014;
    p3_bit_slice_33947 <= p3_bit_slice_33947_comb;
    p3_bit_slice_33948 <= p3_bit_slice_33948_comb;
    p3_bit_slice_33949 <= p3_bit_slice_33949_comb;
    p3_bit_slice_33950 <= p3_bit_slice_33950_comb;
    p3_bit_slice_33951 <= p3_bit_slice_33951_comb;
    p3_bit_slice_33952 <= p3_bit_slice_33952_comb;
    p3_bit_slice_33953 <= p3_bit_slice_33953_comb;
    p3_bit_slice_33954 <= p3_bit_slice_33954_comb;
    p3_array_index_33017 <= p2_array_index_33017;
    p3_array_index_33018 <= p2_array_index_33018;
    p3_array_index_33021 <= p2_array_index_33021;
    p3_array_index_33022 <= p2_array_index_33022;
    p3_bit_slice_34069 <= p3_bit_slice_34069_comb;
    p3_bit_slice_34070 <= p3_bit_slice_34070_comb;
    p3_bit_slice_34071 <= p3_bit_slice_34071_comb;
    p3_bit_slice_34072 <= p3_bit_slice_34072_comb;
    p3_bit_slice_34073 <= p3_bit_slice_34073_comb;
    p3_bit_slice_34074 <= p3_bit_slice_34074_comb;
    p3_bit_slice_34075 <= p3_bit_slice_34075_comb;
    p3_bit_slice_34076 <= p3_bit_slice_34076_comb;
    p3_bit_slice_33029 <= p2_bit_slice_33029;
    p3_bit_slice_33030 <= p2_bit_slice_33030;
    p3_bit_slice_33033 <= p2_bit_slice_33033;
    p3_bit_slice_33034 <= p2_bit_slice_33034;
    p3_umul_33254 <= p2_umul_33254;
    p3_umul_33256 <= p2_umul_33256;
    p3_umul_33267 <= p2_umul_33267;
    p3_umul_33268 <= p2_umul_33268;
    p3_umul_33270 <= p2_umul_33270;
    p3_umul_33272 <= p2_umul_33272;
    p3_umul_33277 <= p2_umul_33277;
    p3_umul_33278 <= p2_umul_33278;
    p3_umul_33286 <= p2_umul_33286;
    p3_umul_33288 <= p2_umul_33288;
    p3_umul_33293 <= p2_umul_33293;
    p3_umul_33294 <= p2_umul_33294;
  end

  // ===== Pipe stage 4:
  wire [31:0] p4_sign_ext_34317_comb;
  wire [31:0] p4_sign_ext_34318_comb;
  wire [31:0] p4_sign_ext_34319_comb;
  wire [31:0] p4_sign_ext_34320_comb;
  wire [31:0] p4_sign_ext_34321_comb;
  wire [31:0] p4_sign_ext_34322_comb;
  wire [31:0] p4_sign_ext_34323_comb;
  wire [31:0] p4_sign_ext_34324_comb;
  wire [31:0] p4_add_34325_comb;
  wire [31:0] p4_add_34327_comb;
  wire [31:0] p4_add_34329_comb;
  wire [31:0] p4_add_34331_comb;
  wire [31:0] p4_umul_34233_comb;
  wire [31:0] p4_umul_34234_comb;
  wire [31:0] p4_umul_34235_comb;
  wire [31:0] p4_umul_34236_comb;
  wire [31:0] p4_umul_34249_comb;
  wire [31:0] p4_umul_34250_comb;
  wire [31:0] p4_umul_34253_comb;
  wire [31:0] p4_umul_34254_comb;
  wire [31:0] p4_umul_34286_comb;
  wire [31:0] p4_umul_34287_comb;
  wire [31:0] p4_umul_34288_comb;
  wire [31:0] p4_umul_34289_comb;
  wire [31:0] p4_sign_ext_34333_comb;
  wire [31:0] p4_sign_ext_34334_comb;
  wire [31:0] p4_sign_ext_34336_comb;
  wire [31:0] p4_sign_ext_34337_comb;
  wire [31:0] p4_sign_ext_34339_comb;
  wire [31:0] p4_sign_ext_34340_comb;
  wire [31:0] p4_sign_ext_34342_comb;
  wire [31:0] p4_sign_ext_34343_comb;
  wire [31:0] p4_umul_34335_comb;
  wire [31:0] p4_umul_34338_comb;
  wire [31:0] p4_umul_34341_comb;
  wire [31:0] p4_umul_34344_comb;
  wire [31:0] p4_umul_34364_comb;
  wire [31:0] p4_umul_34370_comb;
  wire [31:0] p4_umul_34376_comb;
  wire [31:0] p4_umul_34382_comb;
  wire [31:0] p4_umul_34388_comb;
  wire [31:0] p4_umul_34411_comb;
  wire [31:0] p4_add_34270_comb;
  wire [31:0] p4_add_34275_comb;
  wire [31:0] p4_add_34281_comb;
  wire [31:0] p4_add_34294_comb;
  wire [31:0] p4_add_34346_comb;
  wire [31:0] p4_add_34350_comb;
  wire [31:0] p4_add_34354_comb;
  wire [31:0] p4_add_34358_comb;
  wire [31:0] p4_add_34362_comb;
  wire [31:0] p4_add_34391_comb;
  wire [29:0] p4_bit_slice_34348_comb;
  wire [29:0] p4_bit_slice_34352_comb;
  wire [29:0] p4_bit_slice_34356_comb;
  wire [29:0] p4_bit_slice_34360_comb;
  wire [1:0] p4_bit_slice_34368_comb;
  wire [1:0] p4_bit_slice_34374_comb;
  wire [1:0] p4_bit_slice_34380_comb;
  wire [1:0] p4_bit_slice_34386_comb;
  wire [29:0] p4_bit_slice_34393_comb;
  wire [29:0] p4_bit_slice_34397_comb;
  wire [29:0] p4_bit_slice_34401_comb;
  wire [29:0] p4_bit_slice_34405_comb;
  wire [26:0] p4_bit_slice_34410_comb;
  wire [26:0] p4_bit_slice_34415_comb;
  wire [24:0] p4_add_34251_comb;
  wire [24:0] p4_add_34252_comb;
  wire [24:0] p4_add_34255_comb;
  wire [24:0] p4_add_34256_comb;
  wire [24:0] p4_add_34265_comb;
  wire [24:0] p4_add_34266_comb;
  wire [24:0] p4_add_34267_comb;
  wire [24:0] p4_add_34268_comb;
  wire [24:0] p4_add_34311_comb;
  wire [24:0] p4_add_34312_comb;
  wire [24:0] p4_add_34313_comb;
  wire [24:0] p4_add_34314_comb;
  wire [31:0] p4_umul_34272_comb;
  wire [31:0] p4_umul_34273_comb;
  wire [31:0] p4_umul_34284_comb;
  wire [31:0] p4_umul_34285_comb;
  wire [31:0] p4_umul_34290_comb;
  wire [31:0] p4_umul_34291_comb;
  wire [31:0] p4_umul_34305_comb;
  wire [31:0] p4_umul_34306_comb;
  wire [31:0] p4_umul_34307_comb;
  wire [31:0] p4_umul_34308_comb;
  wire [31:0] p4_umul_34315_comb;
  wire [31:0] p4_umul_34316_comb;
  wire [31:0] p4_umul_34365_comb;
  wire [31:0] p4_umul_34371_comb;
  wire [31:0] p4_umul_34377_comb;
  wire [31:0] p4_umul_34383_comb;
  wire [31:0] p4_umul_34389_comb;
  wire [31:0] p4_umul_34394_comb;
  wire [31:0] p4_umul_34395_comb;
  wire [31:0] p4_umul_34396_comb;
  wire [31:0] p4_umul_34398_comb;
  wire [31:0] p4_umul_34399_comb;
  wire [31:0] p4_umul_34400_comb;
  wire [31:0] p4_umul_34402_comb;
  wire [31:0] p4_umul_34403_comb;
  wire [31:0] p4_umul_34404_comb;
  wire [31:0] p4_umul_34406_comb;
  wire [31:0] p4_umul_34407_comb;
  wire [31:0] p4_umul_34408_comb;
  wire [31:0] p4_umul_34412_comb;
  wire [31:0] p4_umul_34413_comb;
  wire [31:0] p4_umul_34416_comb;
  assign p4_sign_ext_34317_comb = {{8{p3_bit_slice_33889[23]}}, p3_bit_slice_33889};
  assign p4_sign_ext_34318_comb = {{8{p3_bit_slice_33890[23]}}, p3_bit_slice_33890};
  assign p4_sign_ext_34319_comb = {{8{p3_bit_slice_33895[23]}}, p3_bit_slice_33895};
  assign p4_sign_ext_34320_comb = {{8{p3_bit_slice_33896[23]}}, p3_bit_slice_33896};
  assign p4_sign_ext_34321_comb = {{8{p3_bit_slice_33901[23]}}, p3_bit_slice_33901};
  assign p4_sign_ext_34322_comb = {{8{p3_bit_slice_33902[23]}}, p3_bit_slice_33902};
  assign p4_sign_ext_34323_comb = {{8{p3_bit_slice_33907[23]}}, p3_bit_slice_33907};
  assign p4_sign_ext_34324_comb = {{8{p3_bit_slice_33908[23]}}, p3_bit_slice_33908};
  assign p4_add_34325_comb = p4_sign_ext_34317_comb + p4_sign_ext_34318_comb;
  assign p4_add_34327_comb = p4_sign_ext_34319_comb + p4_sign_ext_34320_comb;
  assign p4_add_34329_comb = p4_sign_ext_34321_comb + p4_sign_ext_34322_comb;
  assign p4_add_34331_comb = p4_sign_ext_34323_comb + p4_sign_ext_34324_comb;
  assign p4_umul_34233_comb = umul32b_32b_x_8b(p3_sub_33539, 8'hb5);
  assign p4_umul_34234_comb = umul32b_32b_x_8b(p3_sub_33540, 8'hb5);
  assign p4_umul_34235_comb = umul32b_32b_x_8b(p3_sub_33549, 8'hb5);
  assign p4_umul_34236_comb = umul32b_32b_x_8b(p3_sub_33550, 8'hb5);
  assign p4_umul_34249_comb = umul32b_32b_x_8b(p3_sub_33567, 8'hb5);
  assign p4_umul_34250_comb = umul32b_32b_x_8b(p3_sub_33568, 8'hb5);
  assign p4_umul_34253_comb = umul32b_32b_x_8b(p3_sub_33569, 8'hb5);
  assign p4_umul_34254_comb = umul32b_32b_x_8b(p3_sub_33570, 8'hb5);
  assign p4_umul_34286_comb = umul32b_32b_x_8b(p3_sub_33685, 8'hb5);
  assign p4_umul_34287_comb = umul32b_32b_x_8b(p3_sub_33686, 8'hb5);
  assign p4_umul_34288_comb = umul32b_32b_x_8b(p3_sub_33687, 8'hb5);
  assign p4_umul_34289_comb = umul32b_32b_x_8b(p3_sub_33688, 8'hb5);
  assign p4_sign_ext_34333_comb = {{8{p3_bit_slice_33947[23]}}, p3_bit_slice_33947};
  assign p4_sign_ext_34334_comb = {{8{p3_bit_slice_33948[23]}}, p3_bit_slice_33948};
  assign p4_sign_ext_34336_comb = {{8{p3_bit_slice_33949[23]}}, p3_bit_slice_33949};
  assign p4_sign_ext_34337_comb = {{8{p3_bit_slice_33950[23]}}, p3_bit_slice_33950};
  assign p4_sign_ext_34339_comb = {{8{p3_bit_slice_33951[23]}}, p3_bit_slice_33951};
  assign p4_sign_ext_34340_comb = {{8{p3_bit_slice_33952[23]}}, p3_bit_slice_33952};
  assign p4_sign_ext_34342_comb = {{8{p3_bit_slice_33953[23]}}, p3_bit_slice_33953};
  assign p4_sign_ext_34343_comb = {{8{p3_bit_slice_33954[23]}}, p3_bit_slice_33954};
  assign p4_umul_34335_comb = umul32b_32b_x_10b(p4_add_34325_comb, 10'h235);
  assign p4_umul_34338_comb = umul32b_32b_x_10b(p4_add_34327_comb, 10'h235);
  assign p4_umul_34341_comb = umul32b_32b_x_10b(p4_add_34329_comb, 10'h235);
  assign p4_umul_34344_comb = umul32b_32b_x_10b(p4_add_34331_comb, 10'h235);
  assign p4_umul_34364_comb = umul32b_32b_x_12b(p4_sign_ext_34317_comb, 12'h8e4);
  assign p4_umul_34370_comb = umul32b_32b_x_12b(p4_sign_ext_34319_comb, 12'h8e4);
  assign p4_umul_34376_comb = umul32b_32b_x_12b(p4_sign_ext_34321_comb, 12'h8e4);
  assign p4_umul_34382_comb = umul32b_32b_x_12b(p4_sign_ext_34323_comb, 12'h8e4);
  assign p4_umul_34388_comb = umul32b_32b_x_11b(p3_array_index_33017, 11'h620);
  assign p4_umul_34411_comb = umul32b_32b_x_11b(p3_array_index_33021, 11'h620);
  assign p4_add_34270_comb = p3_array_index_32965 + p3_array_index_32966;
  assign p4_add_34275_comb = p3_array_index_32979 + p3_array_index_32980;
  assign p4_add_34281_comb = p3_array_index_32985 + p3_array_index_32986;
  assign p4_add_34294_comb = p3_array_index_32997 + p3_array_index_32998;
  assign p4_add_34346_comb = p4_sign_ext_34333_comb + p4_sign_ext_34334_comb;
  assign p4_add_34350_comb = p4_sign_ext_34336_comb + p4_sign_ext_34337_comb;
  assign p4_add_34354_comb = p4_sign_ext_34339_comb + p4_sign_ext_34340_comb;
  assign p4_add_34358_comb = p4_sign_ext_34342_comb + p4_sign_ext_34343_comb;
  assign p4_add_34362_comb = p3_array_index_33017 + p3_array_index_33018;
  assign p4_add_34391_comb = p3_array_index_33021 + p3_array_index_33022;
  assign p4_bit_slice_34348_comb = p4_umul_34335_comb[31:2];
  assign p4_bit_slice_34352_comb = p4_umul_34338_comb[31:2];
  assign p4_bit_slice_34356_comb = p4_umul_34341_comb[31:2];
  assign p4_bit_slice_34360_comb = p4_umul_34344_comb[31:2];
  assign p4_bit_slice_34368_comb = p4_umul_34335_comb[1:0];
  assign p4_bit_slice_34374_comb = p4_umul_34338_comb[1:0];
  assign p4_bit_slice_34380_comb = p4_umul_34341_comb[1:0];
  assign p4_bit_slice_34386_comb = p4_umul_34344_comb[1:0];
  assign p4_bit_slice_34393_comb = p4_umul_34364_comb[31:2];
  assign p4_bit_slice_34397_comb = p4_umul_34370_comb[31:2];
  assign p4_bit_slice_34401_comb = p4_umul_34376_comb[31:2];
  assign p4_bit_slice_34405_comb = p4_umul_34382_comb[31:2];
  assign p4_bit_slice_34410_comb = p4_umul_34388_comb[31:5];
  assign p4_bit_slice_34415_comb = p4_umul_34411_comb[31:5];
  assign p4_add_34251_comb = p4_umul_34233_comb[31:7] + 25'h000_0001;
  assign p4_add_34252_comb = p4_umul_34234_comb[31:7] + 25'h000_0001;
  assign p4_add_34255_comb = p4_umul_34235_comb[31:7] + 25'h000_0001;
  assign p4_add_34256_comb = p4_umul_34236_comb[31:7] + 25'h000_0001;
  assign p4_add_34265_comb = p4_umul_34249_comb[31:7] + 25'h000_0001;
  assign p4_add_34266_comb = p4_umul_34250_comb[31:7] + 25'h000_0001;
  assign p4_add_34267_comb = p4_umul_34253_comb[31:7] + 25'h000_0001;
  assign p4_add_34268_comb = p4_umul_34254_comb[31:7] + 25'h000_0001;
  assign p4_add_34311_comb = p4_umul_34286_comb[31:7] + 25'h000_0001;
  assign p4_add_34312_comb = p4_umul_34287_comb[31:7] + 25'h000_0001;
  assign p4_add_34313_comb = p4_umul_34288_comb[31:7] + 25'h000_0001;
  assign p4_add_34314_comb = p4_umul_34289_comb[31:7] + 25'h000_0001;
  assign p4_umul_34272_comb = umul32b_32b_x_12b(p3_array_index_32965, 12'h8e4);
  assign p4_umul_34273_comb = umul32b_32b_x_10b(p4_add_34270_comb, 10'h235);
  assign p4_umul_34284_comb = umul32b_32b_x_12b(p3_array_index_32979, 12'h8e4);
  assign p4_umul_34285_comb = umul32b_32b_x_10b(p4_add_34275_comb, 10'h235);
  assign p4_umul_34290_comb = umul32b_32b_x_12b(p4_add_34281_comb, 12'h968);
  assign p4_umul_34291_comb = umul32b_32b_x_12b(p3_array_index_32966, 12'hd4e);
  assign p4_umul_34305_comb = umul32b_32b_x_10b(p3_array_index_32985, 10'h31f);
  assign p4_umul_34306_comb = umul32b_32b_x_12b(p3_array_index_32986, 12'hfb1);
  assign p4_umul_34307_comb = umul32b_32b_x_12b(p4_add_34294_comb, 12'h968);
  assign p4_umul_34308_comb = umul32b_32b_x_12b(p3_array_index_32980, 12'hd4e);
  assign p4_umul_34315_comb = umul32b_32b_x_10b(p3_array_index_32997, 10'h31f);
  assign p4_umul_34316_comb = umul32b_32b_x_12b(p3_array_index_32998, 12'hfb1);
  assign p4_umul_34365_comb = umul32b_32b_x_12b(p4_add_34346_comb, 12'h968);
  assign p4_umul_34371_comb = umul32b_32b_x_12b(p4_add_34350_comb, 12'h968);
  assign p4_umul_34377_comb = umul32b_32b_x_12b(p4_add_34354_comb, 12'h968);
  assign p4_umul_34383_comb = umul32b_32b_x_12b(p4_add_34358_comb, 12'h968);
  assign p4_umul_34389_comb = umul32b_32b_x_11b(p4_add_34362_comb, 11'h454);
  assign p4_umul_34394_comb = umul32b_32b_x_12b(p4_sign_ext_34334_comb, 12'hfb1);
  assign p4_umul_34395_comb = umul32b_32b_x_10b(p4_sign_ext_34333_comb, 10'h31f);
  assign p4_umul_34396_comb = umul32b_32b_x_12b(p4_sign_ext_34318_comb, 12'hd4e);
  assign p4_umul_34398_comb = umul32b_32b_x_12b(p4_sign_ext_34337_comb, 12'hfb1);
  assign p4_umul_34399_comb = umul32b_32b_x_10b(p4_sign_ext_34336_comb, 10'h31f);
  assign p4_umul_34400_comb = umul32b_32b_x_12b(p4_sign_ext_34320_comb, 12'hd4e);
  assign p4_umul_34402_comb = umul32b_32b_x_12b(p4_sign_ext_34340_comb, 12'hfb1);
  assign p4_umul_34403_comb = umul32b_32b_x_10b(p4_sign_ext_34339_comb, 10'h31f);
  assign p4_umul_34404_comb = umul32b_32b_x_12b(p4_sign_ext_34322_comb, 12'hd4e);
  assign p4_umul_34406_comb = umul32b_32b_x_12b(p4_sign_ext_34343_comb, 12'hfb1);
  assign p4_umul_34407_comb = umul32b_32b_x_10b(p4_sign_ext_34342_comb, 10'h31f);
  assign p4_umul_34408_comb = umul32b_32b_x_12b(p4_sign_ext_34324_comb, 12'hd4e);
  assign p4_umul_34412_comb = umul32b_32b_x_11b(p4_add_34391_comb, 11'h454);
  assign p4_umul_34413_comb = umul32b_32b_x_12b(p3_array_index_33018, 12'hec8);
  assign p4_umul_34416_comb = umul32b_32b_x_12b(p3_array_index_33022, 12'hec8);

  // Registers for pipe stage 4:
  reg [20:0] p4_bit_slice_32973;
  reg [20:0] p4_bit_slice_32974;
  reg [20:0] p4_bit_slice_32975;
  reg [20:0] p4_bit_slice_32976;
  reg [20:0] p4_bit_slice_32989;
  reg [20:0] p4_bit_slice_32990;
  reg [20:0] p4_bit_slice_32991;
  reg [20:0] p4_bit_slice_32992;
  reg [20:0] p4_bit_slice_33011;
  reg [20:0] p4_bit_slice_33012;
  reg [20:0] p4_bit_slice_33013;
  reg [20:0] p4_bit_slice_33014;
  reg [29:0] p4_bit_slice_34348;
  reg [29:0] p4_bit_slice_34352;
  reg [29:0] p4_bit_slice_34356;
  reg [29:0] p4_bit_slice_34360;
  reg [1:0] p4_bit_slice_34368;
  reg [1:0] p4_bit_slice_34374;
  reg [1:0] p4_bit_slice_34380;
  reg [1:0] p4_bit_slice_34386;
  reg [29:0] p4_bit_slice_34393;
  reg [29:0] p4_bit_slice_34397;
  reg [29:0] p4_bit_slice_34401;
  reg [29:0] p4_bit_slice_34405;
  reg [26:0] p4_bit_slice_34410;
  reg [23:0] p4_bit_slice_34069;
  reg [23:0] p4_bit_slice_34070;
  reg [23:0] p4_bit_slice_34071;
  reg [23:0] p4_bit_slice_34072;
  reg [23:0] p4_bit_slice_34073;
  reg [23:0] p4_bit_slice_34074;
  reg [23:0] p4_bit_slice_34075;
  reg [23:0] p4_bit_slice_34076;
  reg [20:0] p4_bit_slice_33029;
  reg [20:0] p4_bit_slice_33030;
  reg [26:0] p4_bit_slice_34415;
  reg [20:0] p4_bit_slice_33033;
  reg [20:0] p4_bit_slice_33034;
  reg [24:0] p4_add_34251;
  reg [24:0] p4_add_34252;
  reg [24:0] p4_add_34255;
  reg [24:0] p4_add_34256;
  reg [24:0] p4_add_34265;
  reg [24:0] p4_add_34266;
  reg [24:0] p4_add_34267;
  reg [24:0] p4_add_34268;
  reg [24:0] p4_add_34311;
  reg [24:0] p4_add_34312;
  reg [24:0] p4_add_34313;
  reg [24:0] p4_add_34314;
  reg [31:0] p4_umul_33254;
  reg [31:0] p4_umul_33256;
  reg [31:0] p4_umul_33267;
  reg [31:0] p4_umul_33268;
  reg [31:0] p4_umul_33270;
  reg [31:0] p4_umul_33272;
  reg [31:0] p4_umul_34272;
  reg [31:0] p4_umul_34273;
  reg [31:0] p4_umul_33277;
  reg [31:0] p4_umul_33278;
  reg [31:0] p4_umul_34284;
  reg [31:0] p4_umul_34285;
  reg [31:0] p4_umul_34290;
  reg [31:0] p4_umul_34291;
  reg [31:0] p4_umul_34305;
  reg [31:0] p4_umul_34306;
  reg [31:0] p4_umul_34307;
  reg [31:0] p4_umul_34308;
  reg [31:0] p4_umul_33286;
  reg [31:0] p4_umul_33288;
  reg [31:0] p4_umul_34315;
  reg [31:0] p4_umul_34316;
  reg [31:0] p4_umul_33293;
  reg [31:0] p4_umul_33294;
  reg [31:0] p4_umul_34365;
  reg [31:0] p4_umul_34371;
  reg [31:0] p4_umul_34377;
  reg [31:0] p4_umul_34383;
  reg [31:0] p4_umul_34389;
  reg [31:0] p4_umul_34394;
  reg [31:0] p4_umul_34395;
  reg [31:0] p4_umul_34396;
  reg [31:0] p4_umul_34398;
  reg [31:0] p4_umul_34399;
  reg [31:0] p4_umul_34400;
  reg [31:0] p4_umul_34402;
  reg [31:0] p4_umul_34403;
  reg [31:0] p4_umul_34404;
  reg [31:0] p4_umul_34406;
  reg [31:0] p4_umul_34407;
  reg [31:0] p4_umul_34408;
  reg [31:0] p4_umul_34412;
  reg [31:0] p4_umul_34413;
  reg [31:0] p4_umul_34416;
  always_ff @ (posedge clk) begin
    p4_bit_slice_32973 <= p3_bit_slice_32973;
    p4_bit_slice_32974 <= p3_bit_slice_32974;
    p4_bit_slice_32975 <= p3_bit_slice_32975;
    p4_bit_slice_32976 <= p3_bit_slice_32976;
    p4_bit_slice_32989 <= p3_bit_slice_32989;
    p4_bit_slice_32990 <= p3_bit_slice_32990;
    p4_bit_slice_32991 <= p3_bit_slice_32991;
    p4_bit_slice_32992 <= p3_bit_slice_32992;
    p4_bit_slice_33011 <= p3_bit_slice_33011;
    p4_bit_slice_33012 <= p3_bit_slice_33012;
    p4_bit_slice_33013 <= p3_bit_slice_33013;
    p4_bit_slice_33014 <= p3_bit_slice_33014;
    p4_bit_slice_34348 <= p4_bit_slice_34348_comb;
    p4_bit_slice_34352 <= p4_bit_slice_34352_comb;
    p4_bit_slice_34356 <= p4_bit_slice_34356_comb;
    p4_bit_slice_34360 <= p4_bit_slice_34360_comb;
    p4_bit_slice_34368 <= p4_bit_slice_34368_comb;
    p4_bit_slice_34374 <= p4_bit_slice_34374_comb;
    p4_bit_slice_34380 <= p4_bit_slice_34380_comb;
    p4_bit_slice_34386 <= p4_bit_slice_34386_comb;
    p4_bit_slice_34393 <= p4_bit_slice_34393_comb;
    p4_bit_slice_34397 <= p4_bit_slice_34397_comb;
    p4_bit_slice_34401 <= p4_bit_slice_34401_comb;
    p4_bit_slice_34405 <= p4_bit_slice_34405_comb;
    p4_bit_slice_34410 <= p4_bit_slice_34410_comb;
    p4_bit_slice_34069 <= p3_bit_slice_34069;
    p4_bit_slice_34070 <= p3_bit_slice_34070;
    p4_bit_slice_34071 <= p3_bit_slice_34071;
    p4_bit_slice_34072 <= p3_bit_slice_34072;
    p4_bit_slice_34073 <= p3_bit_slice_34073;
    p4_bit_slice_34074 <= p3_bit_slice_34074;
    p4_bit_slice_34075 <= p3_bit_slice_34075;
    p4_bit_slice_34076 <= p3_bit_slice_34076;
    p4_bit_slice_33029 <= p3_bit_slice_33029;
    p4_bit_slice_33030 <= p3_bit_slice_33030;
    p4_bit_slice_34415 <= p4_bit_slice_34415_comb;
    p4_bit_slice_33033 <= p3_bit_slice_33033;
    p4_bit_slice_33034 <= p3_bit_slice_33034;
    p4_add_34251 <= p4_add_34251_comb;
    p4_add_34252 <= p4_add_34252_comb;
    p4_add_34255 <= p4_add_34255_comb;
    p4_add_34256 <= p4_add_34256_comb;
    p4_add_34265 <= p4_add_34265_comb;
    p4_add_34266 <= p4_add_34266_comb;
    p4_add_34267 <= p4_add_34267_comb;
    p4_add_34268 <= p4_add_34268_comb;
    p4_add_34311 <= p4_add_34311_comb;
    p4_add_34312 <= p4_add_34312_comb;
    p4_add_34313 <= p4_add_34313_comb;
    p4_add_34314 <= p4_add_34314_comb;
    p4_umul_33254 <= p3_umul_33254;
    p4_umul_33256 <= p3_umul_33256;
    p4_umul_33267 <= p3_umul_33267;
    p4_umul_33268 <= p3_umul_33268;
    p4_umul_33270 <= p3_umul_33270;
    p4_umul_33272 <= p3_umul_33272;
    p4_umul_34272 <= p4_umul_34272_comb;
    p4_umul_34273 <= p4_umul_34273_comb;
    p4_umul_33277 <= p3_umul_33277;
    p4_umul_33278 <= p3_umul_33278;
    p4_umul_34284 <= p4_umul_34284_comb;
    p4_umul_34285 <= p4_umul_34285_comb;
    p4_umul_34290 <= p4_umul_34290_comb;
    p4_umul_34291 <= p4_umul_34291_comb;
    p4_umul_34305 <= p4_umul_34305_comb;
    p4_umul_34306 <= p4_umul_34306_comb;
    p4_umul_34307 <= p4_umul_34307_comb;
    p4_umul_34308 <= p4_umul_34308_comb;
    p4_umul_33286 <= p3_umul_33286;
    p4_umul_33288 <= p3_umul_33288;
    p4_umul_34315 <= p4_umul_34315_comb;
    p4_umul_34316 <= p4_umul_34316_comb;
    p4_umul_33293 <= p3_umul_33293;
    p4_umul_33294 <= p3_umul_33294;
    p4_umul_34365 <= p4_umul_34365_comb;
    p4_umul_34371 <= p4_umul_34371_comb;
    p4_umul_34377 <= p4_umul_34377_comb;
    p4_umul_34383 <= p4_umul_34383_comb;
    p4_umul_34389 <= p4_umul_34389_comb;
    p4_umul_34394 <= p4_umul_34394_comb;
    p4_umul_34395 <= p4_umul_34395_comb;
    p4_umul_34396 <= p4_umul_34396_comb;
    p4_umul_34398 <= p4_umul_34398_comb;
    p4_umul_34399 <= p4_umul_34399_comb;
    p4_umul_34400 <= p4_umul_34400_comb;
    p4_umul_34402 <= p4_umul_34402_comb;
    p4_umul_34403 <= p4_umul_34403_comb;
    p4_umul_34404 <= p4_umul_34404_comb;
    p4_umul_34406 <= p4_umul_34406_comb;
    p4_umul_34407 <= p4_umul_34407_comb;
    p4_umul_34408 <= p4_umul_34408_comb;
    p4_umul_34412 <= p4_umul_34412_comb;
    p4_umul_34413 <= p4_umul_34413_comb;
    p4_umul_34416 <= p4_umul_34416_comb;
  end

  // ===== Pipe stage 5:
  wire [23:0] p5_bit_slice_34605_comb;
  wire [23:0] p5_bit_slice_34606_comb;
  wire [23:0] p5_bit_slice_34607_comb;
  wire [23:0] p5_bit_slice_34608_comb;
  wire [23:0] p5_bit_slice_34613_comb;
  wire [23:0] p5_bit_slice_34614_comb;
  wire [23:0] p5_bit_slice_34621_comb;
  wire [23:0] p5_bit_slice_34622_comb;
  wire [23:0] p5_bit_slice_34879_comb;
  wire [23:0] p5_bit_slice_34880_comb;
  wire [23:0] p5_bit_slice_34881_comb;
  wire [23:0] p5_bit_slice_34882_comb;
  wire [31:0] p5_sign_ext_34609_comb;
  wire [31:0] p5_sign_ext_34610_comb;
  wire [31:0] p5_sign_ext_34611_comb;
  wire [31:0] p5_sign_ext_34612_comb;
  wire [31:0] p5_sign_ext_34645_comb;
  wire [31:0] p5_sign_ext_34646_comb;
  wire [31:0] p5_sign_ext_34655_comb;
  wire [31:0] p5_sign_ext_34656_comb;
  wire [31:0] p5_sign_ext_34914_comb;
  wire [31:0] p5_sign_ext_34915_comb;
  wire [31:0] p5_sign_ext_34916_comb;
  wire [31:0] p5_sign_ext_34917_comb;
  wire [29:0] p5_add_34719_comb;
  wire [29:0] p5_add_34790_comb;
  wire [29:0] p5_add_35074_comb;
  wire [29:0] p5_add_35076_comb;
  wire [29:0] p5_add_35078_comb;
  wire [29:0] p5_add_35080_comb;
  wire [26:0] p5_add_35138_comb;
  wire [26:0] p5_add_35178_comb;
  wire [24:0] p5_add_34647_comb;
  wire [20:0] p5_add_34649_comb;
  wire [24:0] p5_add_34651_comb;
  wire [20:0] p5_add_34653_comb;
  wire [24:0] p5_add_34657_comb;
  wire [20:0] p5_add_34659_comb;
  wire [24:0] p5_add_34661_comb;
  wire [20:0] p5_add_34663_comb;
  wire [24:0] p5_add_34665_comb;
  wire [29:0] p5_add_34666_comb;
  wire [24:0] p5_add_34667_comb;
  wire [29:0] p5_add_34668_comb;
  wire [24:0] p5_add_34669_comb;
  wire [28:0] p5_add_34670_comb;
  wire [24:0] p5_add_34671_comb;
  wire [28:0] p5_add_34672_comb;
  wire [24:0] p5_add_34723_comb;
  wire [20:0] p5_add_34725_comb;
  wire [24:0] p5_add_34727_comb;
  wire [20:0] p5_add_34729_comb;
  wire [24:0] p5_add_34739_comb;
  wire [20:0] p5_add_34741_comb;
  wire [24:0] p5_add_34743_comb;
  wire [20:0] p5_add_34745_comb;
  wire [24:0] p5_add_34755_comb;
  wire [29:0] p5_add_34756_comb;
  wire [24:0] p5_add_34757_comb;
  wire [29:0] p5_add_34758_comb;
  wire [24:0] p5_add_34771_comb;
  wire [28:0] p5_add_34772_comb;
  wire [24:0] p5_add_34773_comb;
  wire [28:0] p5_add_34774_comb;
  wire [31:0] p5_concat_34789_comb;
  wire [31:0] p5_concat_34830_comb;
  wire [24:0] p5_add_34981_comb;
  wire [20:0] p5_add_34983_comb;
  wire [24:0] p5_add_34985_comb;
  wire [20:0] p5_add_34987_comb;
  wire [24:0] p5_add_34989_comb;
  wire [20:0] p5_add_34991_comb;
  wire [24:0] p5_add_34993_comb;
  wire [20:0] p5_add_34995_comb;
  wire [24:0] p5_add_34997_comb;
  wire [29:0] p5_add_34998_comb;
  wire [24:0] p5_add_34999_comb;
  wire [29:0] p5_add_35000_comb;
  wire [24:0] p5_add_35001_comb;
  wire [28:0] p5_add_35002_comb;
  wire [24:0] p5_add_35003_comb;
  wire [28:0] p5_add_35004_comb;
  wire [31:0] p5_or_35097_comb;
  wire [31:0] p5_or_35099_comb;
  wire [31:0] p5_or_35101_comb;
  wire [31:0] p5_or_35103_comb;
  wire [20:0] p5_add_35167_comb;
  wire [20:0] p5_add_35213_comb;
  wire [28:0] p5_add_34824_comb;
  wire [31:0] p5_add_34826_comb;
  wire [31:0] p5_add_34827_comb;
  wire [28:0] p5_add_34886_comb;
  wire [31:0] p5_add_34888_comb;
  wire [31:0] p5_add_34889_comb;
  wire [29:0] p5_add_35114_comb;
  wire [31:0] p5_sub_35115_comb;
  wire [31:0] p5_sub_35116_comb;
  wire [31:0] p5_sub_35117_comb;
  wire [29:0] p5_add_35118_comb;
  wire [31:0] p5_sub_35119_comb;
  wire [31:0] p5_sub_35120_comb;
  wire [31:0] p5_sub_35121_comb;
  wire [29:0] p5_add_35122_comb;
  wire [31:0] p5_sub_35123_comb;
  wire [31:0] p5_sub_35124_comb;
  wire [31:0] p5_sub_35125_comb;
  wire [29:0] p5_add_35126_comb;
  wire [31:0] p5_sub_35127_comb;
  wire [31:0] p5_sub_35128_comb;
  wire [31:0] p5_sub_35129_comb;
  wire [24:0] p5_add_35204_comb;
  wire [20:0] p5_add_35206_comb;
  wire [30:0] p5_add_35208_comb;
  wire [24:0] p5_add_35216_comb;
  wire [20:0] p5_add_35218_comb;
  wire [28:0] p5_add_35220_comb;
  wire [24:0] p5_add_35226_comb;
  wire [20:0] p5_add_35228_comb;
  wire [28:0] p5_add_35230_comb;
  wire [24:0] p5_add_35256_comb;
  wire [20:0] p5_add_35258_comb;
  wire [30:0] p5_add_35260_comb;
  wire [24:0] p5_add_35265_comb;
  wire [20:0] p5_add_35267_comb;
  wire [28:0] p5_add_35269_comb;
  wire [24:0] p5_add_35274_comb;
  wire [20:0] p5_add_35276_comb;
  wire [28:0] p5_add_35278_comb;
  wire [29:0] p5_add_34731_comb;
  wire [20:0] p5_add_34733_comb;
  wire [29:0] p5_add_34735_comb;
  wire [20:0] p5_add_34737_comb;
  wire [28:0] p5_add_34747_comb;
  wire [20:0] p5_add_34749_comb;
  wire [28:0] p5_add_34751_comb;
  wire [20:0] p5_add_34753_comb;
  wire [20:0] p5_add_34759_comb;
  wire [20:0] p5_add_34762_comb;
  wire [20:0] p5_add_34765_comb;
  wire [20:0] p5_add_34768_comb;
  wire [20:0] p5_add_34775_comb;
  wire [20:0] p5_add_34778_comb;
  wire [20:0] p5_add_34781_comb;
  wire [20:0] p5_add_34784_comb;
  wire [29:0] p5_add_34831_comb;
  wire [20:0] p5_add_34833_comb;
  wire [29:0] p5_add_34835_comb;
  wire [20:0] p5_add_34837_comb;
  wire [28:0] p5_add_34841_comb;
  wire [20:0] p5_add_34843_comb;
  wire [28:0] p5_add_34845_comb;
  wire [20:0] p5_add_34847_comb;
  wire [20:0] p5_add_34851_comb;
  wire [20:0] p5_add_34854_comb;
  wire [20:0] p5_add_34857_comb;
  wire [20:0] p5_add_34860_comb;
  wire [20:0] p5_add_34865_comb;
  wire [20:0] p5_add_34868_comb;
  wire [20:0] p5_add_34871_comb;
  wire [20:0] p5_add_34874_comb;
  wire [29:0] p5_add_35033_comb;
  wire [20:0] p5_add_35035_comb;
  wire [29:0] p5_add_35037_comb;
  wire [20:0] p5_add_35039_comb;
  wire [28:0] p5_add_35041_comb;
  wire [20:0] p5_add_35043_comb;
  wire [28:0] p5_add_35045_comb;
  wire [20:0] p5_add_35047_comb;
  wire [20:0] p5_add_35049_comb;
  wire [20:0] p5_add_35052_comb;
  wire [20:0] p5_add_35055_comb;
  wire [20:0] p5_add_35058_comb;
  wire [20:0] p5_add_35061_comb;
  wire [20:0] p5_add_35064_comb;
  wire [20:0] p5_add_35067_comb;
  wire [20:0] p5_add_35070_comb;
  wire [28:0] p5_bit_slice_35140_comb;
  wire [28:0] p5_bit_slice_35141_comb;
  wire [28:0] p5_bit_slice_35142_comb;
  wire [28:0] p5_bit_slice_35143_comb;
  wire [28:0] p5_bit_slice_35144_comb;
  wire [28:0] p5_bit_slice_35145_comb;
  wire [28:0] p5_bit_slice_35146_comb;
  wire [28:0] p5_bit_slice_35147_comb;
  wire [28:0] p5_bit_slice_35148_comb;
  wire [28:0] p5_bit_slice_35149_comb;
  wire [28:0] p5_bit_slice_35150_comb;
  wire [28:0] p5_bit_slice_35151_comb;
  wire [28:0] p5_bit_slice_35152_comb;
  wire [28:0] p5_bit_slice_35153_comb;
  wire [28:0] p5_bit_slice_35154_comb;
  wire [28:0] p5_bit_slice_35155_comb;
  wire [31:0] p5_sign_ext_35156_comb;
  wire [31:0] p5_sign_ext_35157_comb;
  wire [31:0] p5_sign_ext_35158_comb;
  wire [31:0] p5_sign_ext_35159_comb;
  wire [31:0] p5_sign_ext_35160_comb;
  wire [31:0] p5_sign_ext_35161_comb;
  wire [31:0] p5_sign_ext_35162_comb;
  wire [31:0] p5_sign_ext_35163_comb;
  wire [31:0] p5_sub_35248_comb;
  wire [29:0] p5_concat_35255_comb;
  wire [31:0] p5_sub_35291_comb;
  wire [29:0] p5_concat_35302_comb;
  wire [28:0] p5_add_34918_comb;
  wire [30:0] p5_add_34920_comb;
  wire [28:0] p5_add_34922_comb;
  wire [28:0] p5_add_34965_comb;
  wire [30:0] p5_add_34969_comb;
  wire [28:0] p5_add_34971_comb;
  wire [31:0] p5_sign_ext_35179_comb;
  wire [31:0] p5_sign_ext_35180_comb;
  wire [31:0] p5_sign_ext_35181_comb;
  wire [31:0] p5_sign_ext_35182_comb;
  wire [31:0] p5_sign_ext_35183_comb;
  wire [31:0] p5_sign_ext_35184_comb;
  wire [31:0] p5_sign_ext_35185_comb;
  wire [31:0] p5_sign_ext_35186_comb;
  wire [31:0] p5_sign_ext_35187_comb;
  wire [31:0] p5_sign_ext_35188_comb;
  wire [31:0] p5_sign_ext_35189_comb;
  wire [31:0] p5_sign_ext_35190_comb;
  wire [31:0] p5_sign_ext_35191_comb;
  wire [31:0] p5_sign_ext_35192_comb;
  wire [31:0] p5_sign_ext_35193_comb;
  wire [31:0] p5_sign_ext_35194_comb;
  wire [31:0] p5_add_35195_comb;
  wire [31:0] p5_add_35197_comb;
  wire [31:0] p5_add_35199_comb;
  wire [31:0] p5_add_35201_comb;
  wire [31:0] p5_add_35288_comb;
  wire [24:0] p5_add_35289_comb;
  wire [28:0] p5_add_35294_comb;
  wire [29:0] p5_add_35296_comb;
  wire [30:0] p5_add_35303_comb;
  wire [29:0] p5_add_35304_comb;
  wire [29:0] p5_add_35308_comb;
  wire [29:0] p5_add_35310_comb;
  wire [31:0] p5_add_35332_comb;
  wire [24:0] p5_add_35333_comb;
  wire [28:0] p5_add_35337_comb;
  wire [29:0] p5_add_35339_comb;
  wire [30:0] p5_add_35344_comb;
  wire [29:0] p5_add_35345_comb;
  wire [29:0] p5_add_35348_comb;
  wire [29:0] p5_add_35350_comb;
  wire [31:0] p5_sub_34839_comb;
  wire [31:0] p5_sub_34840_comb;
  wire [31:0] p5_sub_34849_comb;
  wire [31:0] p5_sub_34850_comb;
  wire [31:0] p5_sub_34863_comb;
  wire [31:0] p5_sub_34864_comb;
  wire [31:0] p5_sub_34877_comb;
  wire [31:0] p5_sub_34878_comb;
  wire [31:0] p5_sub_34927_comb;
  wire [31:0] p5_sub_34928_comb;
  wire [31:0] p5_sub_34929_comb;
  wire [31:0] p5_sub_34930_comb;
  wire [31:0] p5_sub_34931_comb;
  wire [31:0] p5_sub_34932_comb;
  wire [31:0] p5_sub_34933_comb;
  wire [31:0] p5_sub_34934_comb;
  wire [31:0] p5_add_34963_comb;
  wire [31:0] p5_add_35006_comb;
  wire [31:0] p5_sub_35105_comb;
  wire [31:0] p5_sub_35106_comb;
  wire [31:0] p5_sub_35107_comb;
  wire [31:0] p5_sub_35108_comb;
  wire [31:0] p5_sub_35109_comb;
  wire [31:0] p5_sub_35110_comb;
  wire [31:0] p5_sub_35111_comb;
  wire [31:0] p5_sub_35112_comb;
  wire [31:0] p5_add_35236_comb;
  wire [31:0] p5_add_35237_comb;
  wire [31:0] p5_add_35238_comb;
  wire [31:0] p5_add_35239_comb;
  wire [31:0] p5_add_35240_comb;
  wire [31:0] p5_add_35241_comb;
  wire [31:0] p5_add_35242_comb;
  wire [31:0] p5_add_35243_comb;
  wire [31:0] p5_umul_35244_comb;
  wire [31:0] p5_umul_35245_comb;
  wire [31:0] p5_umul_35246_comb;
  wire [31:0] p5_umul_35247_comb;
  wire [31:0] p5_add_35315_comb;
  wire [31:0] p5_add_35316_comb;
  wire [31:0] p5_add_35318_comb;
  wire [31:0] p5_add_35319_comb;
  wire [31:0] p5_add_35321_comb;
  wire [31:0] p5_add_35322_comb;
  wire [31:0] p5_add_35324_comb;
  wire [31:0] p5_add_35325_comb;
  wire [31:0] p5_umul_35359_comb;
  wire [31:0] p5_umul_35360_comb;
  wire [31:0] p5_umul_35361_comb;
  wire [31:0] p5_umul_35362_comb;
  wire [23:0] p5_bit_slice_34894_comb;
  wire [23:0] p5_bit_slice_34895_comb;
  wire [23:0] p5_bit_slice_34900_comb;
  wire [23:0] p5_bit_slice_34901_comb;
  wire [23:0] p5_bit_slice_34906_comb;
  wire [23:0] p5_bit_slice_34907_comb;
  wire [23:0] p5_bit_slice_34912_comb;
  wire [23:0] p5_bit_slice_34913_comb;
  wire [23:0] p5_bit_slice_34973_comb;
  wire [23:0] p5_bit_slice_34974_comb;
  wire [23:0] p5_bit_slice_34975_comb;
  wire [23:0] p5_bit_slice_34976_comb;
  wire [23:0] p5_bit_slice_34977_comb;
  wire [23:0] p5_bit_slice_34978_comb;
  wire [23:0] p5_bit_slice_34979_comb;
  wire [23:0] p5_bit_slice_34980_comb;
  wire [31:0] p5_sub_35005_comb;
  wire [31:0] p5_sub_35008_comb;
  wire [31:0] p5_sub_35027_comb;
  wire [31:0] p5_sub_35028_comb;
  wire [23:0] p5_bit_slice_35130_comb;
  wire [23:0] p5_bit_slice_35131_comb;
  wire [23:0] p5_bit_slice_35132_comb;
  wire [23:0] p5_bit_slice_35133_comb;
  wire [23:0] p5_bit_slice_35134_comb;
  wire [23:0] p5_bit_slice_35135_comb;
  wire [23:0] p5_bit_slice_35136_comb;
  wire [23:0] p5_bit_slice_35137_comb;
  wire [31:0] p5_sub_35280_comb;
  wire [31:0] p5_sub_35281_comb;
  wire [31:0] p5_sub_35282_comb;
  wire [31:0] p5_sub_35283_comb;
  wire [29:0] p5_bit_slice_35284_comb;
  wire [29:0] p5_bit_slice_35285_comb;
  wire [29:0] p5_bit_slice_35286_comb;
  wire [29:0] p5_bit_slice_35287_comb;
  wire [31:0] p5_sub_35352_comb;
  wire [31:0] p5_sub_35354_comb;
  wire [31:0] p5_sub_35356_comb;
  wire [31:0] p5_sub_35358_comb;
  wire [29:0] p5_add_35363_comb;
  wire [31:0] p5_sub_35366_comb;
  wire [31:0] p5_sub_35369_comb;
  wire [31:0] p5_sub_35372_comb;
  wire [26:0] p5_bit_slice_35375_comb;
  wire [26:0] p5_bit_slice_35376_comb;
  wire [26:0] p5_bit_slice_35377_comb;
  wire [26:0] p5_bit_slice_35378_comb;
  wire [29:0] p5_add_35379_comb;
  wire [31:0] p5_sub_35380_comb;
  wire [31:0] p5_sub_35381_comb;
  wire [31:0] p5_sub_35382_comb;
  wire [31:0] p5_add_35383_comb;
  wire [31:0] p5_add_35384_comb;
  wire [31:0] p5_add_35385_comb;
  wire [31:0] p5_add_35386_comb;
  wire [31:0] p5_add_35387_comb;
  wire [31:0] p5_add_35388_comb;
  wire [31:0] p5_add_35389_comb;
  wire [31:0] p5_add_35390_comb;
  wire [31:0] p5_umul_35351_comb;
  wire [31:0] p5_umul_35353_comb;
  wire [31:0] p5_umul_35355_comb;
  wire [31:0] p5_umul_35357_comb;
  assign p5_bit_slice_34605_comb = p4_add_34251[24:1];
  assign p5_bit_slice_34606_comb = p4_add_34252[24:1];
  assign p5_bit_slice_34607_comb = p4_add_34255[24:1];
  assign p5_bit_slice_34608_comb = p4_add_34256[24:1];
  assign p5_bit_slice_34613_comb = p4_add_34265[24:1];
  assign p5_bit_slice_34614_comb = p4_add_34266[24:1];
  assign p5_bit_slice_34621_comb = p4_add_34267[24:1];
  assign p5_bit_slice_34622_comb = p4_add_34268[24:1];
  assign p5_bit_slice_34879_comb = p4_add_34311[24:1];
  assign p5_bit_slice_34880_comb = p4_add_34312[24:1];
  assign p5_bit_slice_34881_comb = p4_add_34313[24:1];
  assign p5_bit_slice_34882_comb = p4_add_34314[24:1];
  assign p5_sign_ext_34609_comb = {{8{p5_bit_slice_34605_comb[23]}}, p5_bit_slice_34605_comb};
  assign p5_sign_ext_34610_comb = {{8{p5_bit_slice_34606_comb[23]}}, p5_bit_slice_34606_comb};
  assign p5_sign_ext_34611_comb = {{8{p5_bit_slice_34607_comb[23]}}, p5_bit_slice_34607_comb};
  assign p5_sign_ext_34612_comb = {{8{p5_bit_slice_34608_comb[23]}}, p5_bit_slice_34608_comb};
  assign p5_sign_ext_34645_comb = {{8{p5_bit_slice_34613_comb[23]}}, p5_bit_slice_34613_comb};
  assign p5_sign_ext_34646_comb = {{8{p5_bit_slice_34614_comb[23]}}, p5_bit_slice_34614_comb};
  assign p5_sign_ext_34655_comb = {{8{p5_bit_slice_34621_comb[23]}}, p5_bit_slice_34621_comb};
  assign p5_sign_ext_34656_comb = {{8{p5_bit_slice_34622_comb[23]}}, p5_bit_slice_34622_comb};
  assign p5_sign_ext_34914_comb = {{8{p5_bit_slice_34879_comb[23]}}, p5_bit_slice_34879_comb};
  assign p5_sign_ext_34915_comb = {{8{p5_bit_slice_34880_comb[23]}}, p5_bit_slice_34880_comb};
  assign p5_sign_ext_34916_comb = {{8{p5_bit_slice_34881_comb[23]}}, p5_bit_slice_34881_comb};
  assign p5_sign_ext_34917_comb = {{8{p5_bit_slice_34882_comb[23]}}, p5_bit_slice_34882_comb};
  assign p5_add_34719_comb = p4_umul_34272[31:2] + p4_umul_34273[31:2];
  assign p5_add_34790_comb = p4_umul_34284[31:2] + p4_umul_34285[31:2];
  assign p5_add_35074_comb = p4_bit_slice_34348 + 30'h0000_0001;
  assign p5_add_35076_comb = p4_bit_slice_34352 + 30'h0000_0001;
  assign p5_add_35078_comb = p4_bit_slice_34356 + 30'h0000_0001;
  assign p5_add_35080_comb = p4_bit_slice_34360 + 30'h0000_0001;
  assign p5_add_35138_comb = p4_bit_slice_34410 + p4_umul_34389[31:5];
  assign p5_add_35178_comb = p4_bit_slice_34415 + p4_umul_34412[31:5];
  assign p5_add_34647_comb = p5_sign_ext_34609_comb[31:7] + 25'h000_0001;
  assign p5_add_34649_comb = p4_umul_33254[31:11] + p4_bit_slice_32974;
  assign p5_add_34651_comb = p5_sign_ext_34610_comb[31:7] + 25'h000_0001;
  assign p5_add_34653_comb = p4_umul_33256[31:11] + p4_bit_slice_32976;
  assign p5_add_34657_comb = p5_sign_ext_34611_comb[31:7] + 25'h000_0001;
  assign p5_add_34659_comb = p4_umul_33267[31:11] + p4_bit_slice_32974;
  assign p5_add_34661_comb = p5_sign_ext_34612_comb[31:7] + 25'h000_0001;
  assign p5_add_34663_comb = p4_umul_33268[31:11] + p4_bit_slice_32976;
  assign p5_add_34665_comb = p4_umul_33267[31:7] + 25'h000_0001;
  assign p5_add_34666_comb = p5_sign_ext_34611_comb[31:2] + p4_umul_33254[31:2];
  assign p5_add_34667_comb = p4_umul_33268[31:7] + 25'h000_0001;
  assign p5_add_34668_comb = p5_sign_ext_34612_comb[31:2] + p4_umul_33256[31:2];
  assign p5_add_34669_comb = p4_umul_33254[31:7] + 25'h000_0001;
  assign p5_add_34670_comb = p5_sign_ext_34609_comb[31:3] + p4_umul_33267[31:3];
  assign p5_add_34671_comb = p4_umul_33256[31:7] + 25'h000_0001;
  assign p5_add_34672_comb = p5_sign_ext_34610_comb[31:3] + p4_umul_33268[31:3];
  assign p5_add_34723_comb = p5_sign_ext_34645_comb[31:7] + 25'h000_0001;
  assign p5_add_34725_comb = p4_umul_33270[31:11] + p4_bit_slice_32990;
  assign p5_add_34727_comb = p5_sign_ext_34646_comb[31:7] + 25'h000_0001;
  assign p5_add_34729_comb = p4_umul_33272[31:11] + p4_bit_slice_32992;
  assign p5_add_34739_comb = p5_sign_ext_34655_comb[31:7] + 25'h000_0001;
  assign p5_add_34741_comb = p4_umul_33277[31:11] + p4_bit_slice_32990;
  assign p5_add_34743_comb = p5_sign_ext_34656_comb[31:7] + 25'h000_0001;
  assign p5_add_34745_comb = p4_umul_33278[31:11] + p4_bit_slice_32992;
  assign p5_add_34755_comb = p4_umul_33277[31:7] + 25'h000_0001;
  assign p5_add_34756_comb = p5_sign_ext_34655_comb[31:2] + p4_umul_33270[31:2];
  assign p5_add_34757_comb = p4_umul_33278[31:7] + 25'h000_0001;
  assign p5_add_34758_comb = p5_sign_ext_34656_comb[31:2] + p4_umul_33272[31:2];
  assign p5_add_34771_comb = p4_umul_33270[31:7] + 25'h000_0001;
  assign p5_add_34772_comb = p5_sign_ext_34645_comb[31:3] + p4_umul_33277[31:3];
  assign p5_add_34773_comb = p4_umul_33272[31:7] + 25'h000_0001;
  assign p5_add_34774_comb = p5_sign_ext_34646_comb[31:3] + p4_umul_33278[31:3];
  assign p5_concat_34789_comb = {p5_add_34719_comb, p4_umul_34273[1:0]};
  assign p5_concat_34830_comb = {p5_add_34790_comb, p4_umul_34285[1:0]};
  assign p5_add_34981_comb = p5_sign_ext_34914_comb[31:7] + 25'h000_0001;
  assign p5_add_34983_comb = p4_umul_33286[31:11] + p4_bit_slice_33012;
  assign p5_add_34985_comb = p5_sign_ext_34915_comb[31:7] + 25'h000_0001;
  assign p5_add_34987_comb = p4_umul_33288[31:11] + p4_bit_slice_33014;
  assign p5_add_34989_comb = p5_sign_ext_34916_comb[31:7] + 25'h000_0001;
  assign p5_add_34991_comb = p4_umul_33293[31:11] + p4_bit_slice_33012;
  assign p5_add_34993_comb = p5_sign_ext_34917_comb[31:7] + 25'h000_0001;
  assign p5_add_34995_comb = p4_umul_33294[31:11] + p4_bit_slice_33014;
  assign p5_add_34997_comb = p4_umul_33293[31:7] + 25'h000_0001;
  assign p5_add_34998_comb = p5_sign_ext_34916_comb[31:2] + p4_umul_33286[31:2];
  assign p5_add_34999_comb = p4_umul_33294[31:7] + 25'h000_0001;
  assign p5_add_35000_comb = p5_sign_ext_34917_comb[31:2] + p4_umul_33288[31:2];
  assign p5_add_35001_comb = p4_umul_33286[31:7] + 25'h000_0001;
  assign p5_add_35002_comb = p5_sign_ext_34914_comb[31:3] + p4_umul_33293[31:3];
  assign p5_add_35003_comb = p4_umul_33288[31:7] + 25'h000_0001;
  assign p5_add_35004_comb = p5_sign_ext_34915_comb[31:3] + p4_umul_33294[31:3];
  assign p5_or_35097_comb = p4_umul_34365 | 32'h0000_0004;
  assign p5_or_35099_comb = p4_umul_34371 | 32'h0000_0004;
  assign p5_or_35101_comb = p4_umul_34377 | 32'h0000_0004;
  assign p5_or_35103_comb = p4_umul_34383 | 32'h0000_0004;
  assign p5_add_35167_comb = p4_bit_slice_33029 + p4_bit_slice_33030;
  assign p5_add_35213_comb = p4_bit_slice_33033 + p4_bit_slice_33034;
  assign p5_add_34824_comb = p4_umul_34290[31:3] + p4_umul_34291[31:3];
  assign p5_add_34826_comb = p4_umul_34305 + p5_concat_34789_comb;
  assign p5_add_34827_comb = p4_umul_34306 + p4_umul_34273;
  assign p5_add_34886_comb = p4_umul_34307[31:3] + p4_umul_34308[31:3];
  assign p5_add_34888_comb = p4_umul_34315 + p5_concat_34830_comb;
  assign p5_add_34889_comb = p4_umul_34316 + p4_umul_34285;
  assign p5_add_35114_comb = p4_bit_slice_34393 + p5_add_35074_comb;
  assign p5_sub_35115_comb = p5_or_35097_comb - p4_umul_34394;
  assign p5_sub_35116_comb = p5_or_35097_comb - p4_umul_34395;
  assign p5_sub_35117_comb = {p5_add_35074_comb, p4_bit_slice_34368} - p4_umul_34396;
  assign p5_add_35118_comb = p4_bit_slice_34397 + p5_add_35076_comb;
  assign p5_sub_35119_comb = p5_or_35099_comb - p4_umul_34398;
  assign p5_sub_35120_comb = p5_or_35099_comb - p4_umul_34399;
  assign p5_sub_35121_comb = {p5_add_35076_comb, p4_bit_slice_34374} - p4_umul_34400;
  assign p5_add_35122_comb = p4_bit_slice_34401 + p5_add_35078_comb;
  assign p5_sub_35123_comb = p5_or_35101_comb - p4_umul_34402;
  assign p5_sub_35124_comb = p5_or_35101_comb - p4_umul_34403;
  assign p5_sub_35125_comb = {p5_add_35078_comb, p4_bit_slice_34380} - p4_umul_34404;
  assign p5_add_35126_comb = p4_bit_slice_34405 + p5_add_35080_comb;
  assign p5_sub_35127_comb = p5_or_35103_comb - p4_umul_34406;
  assign p5_sub_35128_comb = p5_or_35103_comb - p4_umul_34407;
  assign p5_sub_35129_comb = {p5_add_35080_comb, p4_bit_slice_34386} - p4_umul_34408;
  assign p5_add_35204_comb = p4_umul_34290[31:7] + 25'h000_0001;
  assign p5_add_35206_comb = p4_umul_34273[31:11] + p5_add_35167_comb;
  assign p5_add_35208_comb = p4_umul_34306[31:1] + p4_umul_34291[31:1];
  assign p5_add_35216_comb = p4_umul_34306[31:7] + 25'h000_0001;
  assign p5_add_35218_comb = p4_umul_34291[31:11] + p5_add_35167_comb;
  assign p5_add_35220_comb = p4_umul_34290[31:3] + p4_umul_34273[31:3];
  assign p5_add_35226_comb = p4_umul_34305[31:7] + 25'h000_0001;
  assign p5_add_35228_comb = p5_add_35138_comb[26:6] + p5_add_35167_comb;
  assign p5_add_35230_comb = p4_umul_34290[31:3] + p4_umul_34272[31:3];
  assign p5_add_35256_comb = p4_umul_34307[31:7] + 25'h000_0001;
  assign p5_add_35258_comb = p4_umul_34285[31:11] + p5_add_35213_comb;
  assign p5_add_35260_comb = p4_umul_34316[31:1] + p4_umul_34308[31:1];
  assign p5_add_35265_comb = p4_umul_34316[31:7] + 25'h000_0001;
  assign p5_add_35267_comb = p4_umul_34308[31:11] + p5_add_35213_comb;
  assign p5_add_35269_comb = p4_umul_34307[31:3] + p4_umul_34285[31:3];
  assign p5_add_35274_comb = p4_umul_34315[31:7] + 25'h000_0001;
  assign p5_add_35276_comb = p5_add_35178_comb[26:6] + p5_add_35213_comb;
  assign p5_add_35278_comb = p4_umul_34307[31:3] + p4_umul_34284[31:3];
  assign p5_add_34731_comb = {p5_add_34647_comb, p4_add_34251[7:3]} + {p5_add_34649_comb, p4_umul_33254[10:2]};
  assign p5_add_34733_comb = p4_umul_33267[31:11] + p4_bit_slice_32973;
  assign p5_add_34735_comb = {p5_add_34651_comb, p4_add_34252[7:3]} + {p5_add_34653_comb, p4_umul_33256[10:2]};
  assign p5_add_34737_comb = p4_umul_33268[31:11] + p4_bit_slice_32975;
  assign p5_add_34747_comb = {p5_add_34657_comb, p4_add_34255[7:4]} + {p5_add_34659_comb, p4_umul_33267[10:3]};
  assign p5_add_34749_comb = p4_umul_33254[31:11] + p4_bit_slice_32973;
  assign p5_add_34751_comb = {p5_add_34661_comb, p4_add_34256[7:4]} + {p5_add_34663_comb, p4_umul_33268[10:3]};
  assign p5_add_34753_comb = p4_umul_33256[31:11] + p4_bit_slice_32975;
  assign p5_add_34759_comb = p5_add_34665_comb[24:4] + p4_bit_slice_32974;
  assign p5_add_34762_comb = p5_add_34666_comb[29:9] + p4_bit_slice_32973;
  assign p5_add_34765_comb = p5_add_34667_comb[24:4] + p4_bit_slice_32976;
  assign p5_add_34768_comb = p5_add_34668_comb[29:9] + p4_bit_slice_32975;
  assign p5_add_34775_comb = p5_add_34669_comb[24:4] + p4_bit_slice_32974;
  assign p5_add_34778_comb = p5_add_34670_comb[28:8] + p4_bit_slice_32973;
  assign p5_add_34781_comb = p5_add_34671_comb[24:4] + p4_bit_slice_32976;
  assign p5_add_34784_comb = p5_add_34672_comb[28:8] + p4_bit_slice_32975;
  assign p5_add_34831_comb = {p5_add_34723_comb, p4_add_34265[7:3]} + {p5_add_34725_comb, p4_umul_33270[10:2]};
  assign p5_add_34833_comb = p4_umul_33277[31:11] + p4_bit_slice_32989;
  assign p5_add_34835_comb = {p5_add_34727_comb, p4_add_34266[7:3]} + {p5_add_34729_comb, p4_umul_33272[10:2]};
  assign p5_add_34837_comb = p4_umul_33278[31:11] + p4_bit_slice_32991;
  assign p5_add_34841_comb = {p5_add_34739_comb, p4_add_34267[7:4]} + {p5_add_34741_comb, p4_umul_33277[10:3]};
  assign p5_add_34843_comb = p4_umul_33270[31:11] + p4_bit_slice_32989;
  assign p5_add_34845_comb = {p5_add_34743_comb, p4_add_34268[7:4]} + {p5_add_34745_comb, p4_umul_33278[10:3]};
  assign p5_add_34847_comb = p4_umul_33272[31:11] + p4_bit_slice_32991;
  assign p5_add_34851_comb = p5_add_34755_comb[24:4] + p4_bit_slice_32990;
  assign p5_add_34854_comb = p5_add_34756_comb[29:9] + p4_bit_slice_32989;
  assign p5_add_34857_comb = p5_add_34757_comb[24:4] + p4_bit_slice_32992;
  assign p5_add_34860_comb = p5_add_34758_comb[29:9] + p4_bit_slice_32991;
  assign p5_add_34865_comb = p5_add_34771_comb[24:4] + p4_bit_slice_32990;
  assign p5_add_34868_comb = p5_add_34772_comb[28:8] + p4_bit_slice_32989;
  assign p5_add_34871_comb = p5_add_34773_comb[24:4] + p4_bit_slice_32992;
  assign p5_add_34874_comb = p5_add_34774_comb[28:8] + p4_bit_slice_32991;
  assign p5_add_35033_comb = {p5_add_34981_comb, p4_add_34311[7:3]} + {p5_add_34983_comb, p4_umul_33286[10:2]};
  assign p5_add_35035_comb = p4_umul_33293[31:11] + p4_bit_slice_33011;
  assign p5_add_35037_comb = {p5_add_34985_comb, p4_add_34312[7:3]} + {p5_add_34987_comb, p4_umul_33288[10:2]};
  assign p5_add_35039_comb = p4_umul_33294[31:11] + p4_bit_slice_33013;
  assign p5_add_35041_comb = {p5_add_34989_comb, p4_add_34313[7:4]} + {p5_add_34991_comb, p4_umul_33293[10:3]};
  assign p5_add_35043_comb = p4_umul_33286[31:11] + p4_bit_slice_33011;
  assign p5_add_35045_comb = {p5_add_34993_comb, p4_add_34314[7:4]} + {p5_add_34995_comb, p4_umul_33294[10:3]};
  assign p5_add_35047_comb = p4_umul_33288[31:11] + p4_bit_slice_33013;
  assign p5_add_35049_comb = p5_add_34997_comb[24:4] + p4_bit_slice_33012;
  assign p5_add_35052_comb = p5_add_34998_comb[29:9] + p4_bit_slice_33011;
  assign p5_add_35055_comb = p5_add_34999_comb[24:4] + p4_bit_slice_33014;
  assign p5_add_35058_comb = p5_add_35000_comb[29:9] + p4_bit_slice_33013;
  assign p5_add_35061_comb = p5_add_35001_comb[24:4] + p4_bit_slice_33012;
  assign p5_add_35064_comb = p5_add_35002_comb[28:8] + p4_bit_slice_33011;
  assign p5_add_35067_comb = p5_add_35003_comb[24:4] + p4_bit_slice_33014;
  assign p5_add_35070_comb = p5_add_35004_comb[28:8] + p4_bit_slice_33013;
  assign p5_bit_slice_35140_comb = p5_add_35114_comb[29:1];
  assign p5_bit_slice_35141_comb = p5_sub_35115_comb[31:3];
  assign p5_bit_slice_35142_comb = p5_sub_35116_comb[31:3];
  assign p5_bit_slice_35143_comb = p5_sub_35117_comb[31:3];
  assign p5_bit_slice_35144_comb = p5_add_35118_comb[29:1];
  assign p5_bit_slice_35145_comb = p5_sub_35119_comb[31:3];
  assign p5_bit_slice_35146_comb = p5_sub_35120_comb[31:3];
  assign p5_bit_slice_35147_comb = p5_sub_35121_comb[31:3];
  assign p5_bit_slice_35148_comb = p5_add_35122_comb[29:1];
  assign p5_bit_slice_35149_comb = p5_sub_35123_comb[31:3];
  assign p5_bit_slice_35150_comb = p5_sub_35124_comb[31:3];
  assign p5_bit_slice_35151_comb = p5_sub_35125_comb[31:3];
  assign p5_bit_slice_35152_comb = p5_add_35126_comb[29:1];
  assign p5_bit_slice_35153_comb = p5_sub_35127_comb[31:3];
  assign p5_bit_slice_35154_comb = p5_sub_35128_comb[31:3];
  assign p5_bit_slice_35155_comb = p5_sub_35129_comb[31:3];
  assign p5_sign_ext_35156_comb = {{8{p4_bit_slice_34069[23]}}, p4_bit_slice_34069};
  assign p5_sign_ext_35157_comb = {{8{p4_bit_slice_34070[23]}}, p4_bit_slice_34070};
  assign p5_sign_ext_35158_comb = {{8{p4_bit_slice_34071[23]}}, p4_bit_slice_34071};
  assign p5_sign_ext_35159_comb = {{8{p4_bit_slice_34072[23]}}, p4_bit_slice_34072};
  assign p5_sign_ext_35160_comb = {{8{p4_bit_slice_34073[23]}}, p4_bit_slice_34073};
  assign p5_sign_ext_35161_comb = {{8{p4_bit_slice_34074[23]}}, p4_bit_slice_34074};
  assign p5_sign_ext_35162_comb = {{8{p4_bit_slice_34075[23]}}, p4_bit_slice_34075};
  assign p5_sign_ext_35163_comb = {{8{p4_bit_slice_34076[23]}}, p4_bit_slice_34076};
  assign p5_sub_35248_comb = p4_umul_34290 - p4_umul_34305;
  assign p5_concat_35255_comb = {p5_add_35138_comb, p4_umul_34389[4:2]};
  assign p5_sub_35291_comb = p4_umul_34307 - p4_umul_34315;
  assign p5_concat_35302_comb = {p5_add_35178_comb, p4_umul_34412[4:2]};
  assign p5_add_34918_comb = p5_add_34824_comb + p4_umul_34290[31:3];
  assign p5_add_34920_comb = {p5_add_34824_comb, p4_umul_34291[2:1]} + p5_add_34826_comb[31:1];
  assign p5_add_34922_comb = p5_add_34827_comb[31:3] + p4_umul_34290[31:3];
  assign p5_add_34965_comb = p5_add_34886_comb + p4_umul_34307[31:3];
  assign p5_add_34969_comb = {p5_add_34886_comb, p4_umul_34308[2:1]} + p5_add_34888_comb[31:1];
  assign p5_add_34971_comb = p5_add_34889_comb[31:3] + p4_umul_34307[31:3];
  assign p5_sign_ext_35179_comb = {{3{p5_bit_slice_35140_comb[28]}}, p5_bit_slice_35140_comb};
  assign p5_sign_ext_35180_comb = {{3{p5_bit_slice_35141_comb[28]}}, p5_bit_slice_35141_comb};
  assign p5_sign_ext_35181_comb = {{3{p5_bit_slice_35142_comb[28]}}, p5_bit_slice_35142_comb};
  assign p5_sign_ext_35182_comb = {{3{p5_bit_slice_35143_comb[28]}}, p5_bit_slice_35143_comb};
  assign p5_sign_ext_35183_comb = {{3{p5_bit_slice_35144_comb[28]}}, p5_bit_slice_35144_comb};
  assign p5_sign_ext_35184_comb = {{3{p5_bit_slice_35145_comb[28]}}, p5_bit_slice_35145_comb};
  assign p5_sign_ext_35185_comb = {{3{p5_bit_slice_35146_comb[28]}}, p5_bit_slice_35146_comb};
  assign p5_sign_ext_35186_comb = {{3{p5_bit_slice_35147_comb[28]}}, p5_bit_slice_35147_comb};
  assign p5_sign_ext_35187_comb = {{3{p5_bit_slice_35148_comb[28]}}, p5_bit_slice_35148_comb};
  assign p5_sign_ext_35188_comb = {{3{p5_bit_slice_35149_comb[28]}}, p5_bit_slice_35149_comb};
  assign p5_sign_ext_35189_comb = {{3{p5_bit_slice_35150_comb[28]}}, p5_bit_slice_35150_comb};
  assign p5_sign_ext_35190_comb = {{3{p5_bit_slice_35151_comb[28]}}, p5_bit_slice_35151_comb};
  assign p5_sign_ext_35191_comb = {{3{p5_bit_slice_35152_comb[28]}}, p5_bit_slice_35152_comb};
  assign p5_sign_ext_35192_comb = {{3{p5_bit_slice_35153_comb[28]}}, p5_bit_slice_35153_comb};
  assign p5_sign_ext_35193_comb = {{3{p5_bit_slice_35154_comb[28]}}, p5_bit_slice_35154_comb};
  assign p5_sign_ext_35194_comb = {{3{p5_bit_slice_35155_comb[28]}}, p5_bit_slice_35155_comb};
  assign p5_add_35195_comb = p5_sign_ext_35156_comb + p5_sign_ext_35157_comb;
  assign p5_add_35197_comb = p5_sign_ext_35158_comb + p5_sign_ext_35159_comb;
  assign p5_add_35199_comb = p5_sign_ext_35160_comb + p5_sign_ext_35161_comb;
  assign p5_add_35201_comb = p5_sign_ext_35162_comb + p5_sign_ext_35163_comb;
  assign p5_add_35288_comb = p5_sub_35248_comb + p5_concat_34789_comb;
  assign p5_add_35289_comb = p5_add_35138_comb[26:2] + {p5_add_35167_comb, 4'h1};
  assign p5_add_35294_comb = {p5_add_35204_comb, p4_umul_34290[6:3]} + {p5_add_35206_comb, p4_umul_34273[10:3]};
  assign p5_add_35296_comb = p5_add_35208_comb[30:1] + p5_concat_35255_comb;
  assign p5_add_35303_comb = {p5_add_35216_comb, p4_umul_34306[6:1]} + {p5_add_35218_comb, p4_umul_34291[10:1]};
  assign p5_add_35304_comb = {p5_add_35220_comb, p4_umul_34273[2]} + p5_concat_35255_comb;
  assign p5_add_35308_comb = {p5_add_35226_comb, p4_umul_34305[6:2]} + {p5_add_35228_comb, p5_add_35138_comb[5:0], p4_umul_34389[4:2]};
  assign p5_add_35310_comb = {p5_add_35230_comb, p4_umul_34272[2]} + p4_umul_34273[31:2];
  assign p5_add_35332_comb = p5_sub_35291_comb + p5_concat_34830_comb;
  assign p5_add_35333_comb = p5_add_35178_comb[26:2] + {p5_add_35213_comb, 4'h1};
  assign p5_add_35337_comb = {p5_add_35256_comb, p4_umul_34307[6:3]} + {p5_add_35258_comb, p4_umul_34285[10:3]};
  assign p5_add_35339_comb = p5_add_35260_comb[30:1] + p5_concat_35302_comb;
  assign p5_add_35344_comb = {p5_add_35265_comb, p4_umul_34316[6:1]} + {p5_add_35267_comb, p4_umul_34308[10:1]};
  assign p5_add_35345_comb = {p5_add_35269_comb, p4_umul_34285[2]} + p5_concat_35302_comb;
  assign p5_add_35348_comb = {p5_add_35274_comb, p4_umul_34315[6:2]} + {p5_add_35276_comb, p5_add_35178_comb[5:0], p4_umul_34412[4:2]};
  assign p5_add_35350_comb = {p5_add_35278_comb, p4_umul_34284[2]} + p4_umul_34285[31:2];
  assign p5_sub_34839_comb = {p5_add_34731_comb, p4_add_34251[2:1]} - {p5_add_34733_comb, p4_umul_33267[10:0]};
  assign p5_sub_34840_comb = {p5_add_34735_comb, p4_add_34252[2:1]} - {p5_add_34737_comb, p4_umul_33268[10:0]};
  assign p5_sub_34849_comb = {p5_add_34747_comb, p4_add_34255[3:1]} - {p5_add_34749_comb, p4_umul_33254[10:0]};
  assign p5_sub_34850_comb = {p5_add_34751_comb, p4_add_34256[3:1]} - {p5_add_34753_comb, p4_umul_33256[10:0]};
  assign p5_sub_34863_comb = {p5_add_34759_comb, p5_add_34665_comb[3:0], p4_umul_33267[6:0]} - {p5_add_34762_comb, p5_add_34666_comb[8:0], p4_add_34255[2:1]};
  assign p5_sub_34864_comb = {p5_add_34765_comb, p5_add_34667_comb[3:0], p4_umul_33268[6:0]} - {p5_add_34768_comb, p5_add_34668_comb[8:0], p4_add_34256[2:1]};
  assign p5_sub_34877_comb = {p5_add_34775_comb, p5_add_34669_comb[3:0], p4_umul_33254[6:0]} - {p5_add_34778_comb, p5_add_34670_comb[7:0], p4_add_34251[3:1]};
  assign p5_sub_34878_comb = {p5_add_34781_comb, p5_add_34671_comb[3:0], p4_umul_33256[6:0]} - {p5_add_34784_comb, p5_add_34672_comb[7:0], p4_add_34252[3:1]};
  assign p5_sub_34927_comb = {p5_add_34831_comb, p4_add_34265[2:1]} - {p5_add_34833_comb, p4_umul_33277[10:0]};
  assign p5_sub_34928_comb = {p5_add_34835_comb, p4_add_34266[2:1]} - {p5_add_34837_comb, p4_umul_33278[10:0]};
  assign p5_sub_34929_comb = {p5_add_34841_comb, p4_add_34267[3:1]} - {p5_add_34843_comb, p4_umul_33270[10:0]};
  assign p5_sub_34930_comb = {p5_add_34845_comb, p4_add_34268[3:1]} - {p5_add_34847_comb, p4_umul_33272[10:0]};
  assign p5_sub_34931_comb = {p5_add_34851_comb, p5_add_34755_comb[3:0], p4_umul_33277[6:0]} - {p5_add_34854_comb, p5_add_34756_comb[8:0], p4_add_34267[2:1]};
  assign p5_sub_34932_comb = {p5_add_34857_comb, p5_add_34757_comb[3:0], p4_umul_33278[6:0]} - {p5_add_34860_comb, p5_add_34758_comb[8:0], p4_add_34268[2:1]};
  assign p5_sub_34933_comb = {p5_add_34865_comb, p5_add_34771_comb[3:0], p4_umul_33270[6:0]} - {p5_add_34868_comb, p5_add_34772_comb[7:0], p4_add_34265[3:1]};
  assign p5_sub_34934_comb = {p5_add_34871_comb, p5_add_34773_comb[3:0], p4_umul_33272[6:0]} - {p5_add_34874_comb, p5_add_34774_comb[7:0], p4_add_34266[3:1]};
  assign p5_add_34963_comb = p5_add_34826_comb + p5_add_34827_comb;
  assign p5_add_35006_comb = p5_add_34888_comb + p5_add_34889_comb;
  assign p5_sub_35105_comb = {p5_add_35033_comb, p4_add_34311[2:1]} - {p5_add_35035_comb, p4_umul_33293[10:0]};
  assign p5_sub_35106_comb = {p5_add_35037_comb, p4_add_34312[2:1]} - {p5_add_35039_comb, p4_umul_33294[10:0]};
  assign p5_sub_35107_comb = {p5_add_35041_comb, p4_add_34313[3:1]} - {p5_add_35043_comb, p4_umul_33286[10:0]};
  assign p5_sub_35108_comb = {p5_add_35045_comb, p4_add_34314[3:1]} - {p5_add_35047_comb, p4_umul_33288[10:0]};
  assign p5_sub_35109_comb = {p5_add_35049_comb, p5_add_34997_comb[3:0], p4_umul_33293[6:0]} - {p5_add_35052_comb, p5_add_34998_comb[8:0], p4_add_34313[2:1]};
  assign p5_sub_35110_comb = {p5_add_35055_comb, p5_add_34999_comb[3:0], p4_umul_33294[6:0]} - {p5_add_35058_comb, p5_add_35000_comb[8:0], p4_add_34314[2:1]};
  assign p5_sub_35111_comb = {p5_add_35061_comb, p5_add_35001_comb[3:0], p4_umul_33286[6:0]} - {p5_add_35064_comb, p5_add_35002_comb[7:0], p4_add_34311[3:1]};
  assign p5_sub_35112_comb = {p5_add_35067_comb, p5_add_35003_comb[3:0], p4_umul_33288[6:0]} - {p5_add_35070_comb, p5_add_35004_comb[7:0], p4_add_34312[3:1]};
  assign p5_add_35236_comb = p5_sign_ext_35179_comb + p5_sign_ext_35180_comb;
  assign p5_add_35237_comb = p5_sign_ext_35181_comb + p5_sign_ext_35182_comb;
  assign p5_add_35238_comb = p5_sign_ext_35183_comb + p5_sign_ext_35184_comb;
  assign p5_add_35239_comb = p5_sign_ext_35185_comb + p5_sign_ext_35186_comb;
  assign p5_add_35240_comb = p5_sign_ext_35187_comb + p5_sign_ext_35188_comb;
  assign p5_add_35241_comb = p5_sign_ext_35189_comb + p5_sign_ext_35190_comb;
  assign p5_add_35242_comb = p5_sign_ext_35191_comb + p5_sign_ext_35192_comb;
  assign p5_add_35243_comb = p5_sign_ext_35193_comb + p5_sign_ext_35194_comb;
  assign p5_umul_35244_comb = umul32b_32b_x_11b(p5_add_35195_comb, 11'h454);
  assign p5_umul_35245_comb = umul32b_32b_x_11b(p5_add_35197_comb, 11'h454);
  assign p5_umul_35246_comb = umul32b_32b_x_11b(p5_add_35199_comb, 11'h454);
  assign p5_umul_35247_comb = umul32b_32b_x_11b(p5_add_35201_comb, 11'h454);
  assign p5_add_35315_comb = p5_sign_ext_35179_comb + p5_sign_ext_35182_comb;
  assign p5_add_35316_comb = p5_sign_ext_35181_comb + p5_sign_ext_35180_comb;
  assign p5_add_35318_comb = p5_sign_ext_35183_comb + p5_sign_ext_35186_comb;
  assign p5_add_35319_comb = p5_sign_ext_35185_comb + p5_sign_ext_35184_comb;
  assign p5_add_35321_comb = p5_sign_ext_35187_comb + p5_sign_ext_35190_comb;
  assign p5_add_35322_comb = p5_sign_ext_35189_comb + p5_sign_ext_35188_comb;
  assign p5_add_35324_comb = p5_sign_ext_35191_comb + p5_sign_ext_35194_comb;
  assign p5_add_35325_comb = p5_sign_ext_35193_comb + p5_sign_ext_35192_comb;
  assign p5_umul_35359_comb = umul32b_32b_x_11b(p5_sign_ext_35156_comb, 11'h620);
  assign p5_umul_35360_comb = umul32b_32b_x_11b(p5_sign_ext_35158_comb, 11'h620);
  assign p5_umul_35361_comb = umul32b_32b_x_11b(p5_sign_ext_35160_comb, 11'h620);
  assign p5_umul_35362_comb = umul32b_32b_x_11b(p5_sign_ext_35162_comb, 11'h620);
  assign p5_bit_slice_34894_comb = p5_sub_34839_comb[31:8];
  assign p5_bit_slice_34895_comb = p5_sub_34840_comb[31:8];
  assign p5_bit_slice_34900_comb = p5_sub_34849_comb[31:8];
  assign p5_bit_slice_34901_comb = p5_sub_34850_comb[31:8];
  assign p5_bit_slice_34906_comb = p5_sub_34863_comb[31:8];
  assign p5_bit_slice_34907_comb = p5_sub_34864_comb[31:8];
  assign p5_bit_slice_34912_comb = p5_sub_34877_comb[31:8];
  assign p5_bit_slice_34913_comb = p5_sub_34878_comb[31:8];
  assign p5_bit_slice_34973_comb = p5_sub_34927_comb[31:8];
  assign p5_bit_slice_34974_comb = p5_sub_34928_comb[31:8];
  assign p5_bit_slice_34975_comb = p5_sub_34929_comb[31:8];
  assign p5_bit_slice_34976_comb = p5_sub_34930_comb[31:8];
  assign p5_bit_slice_34977_comb = p5_sub_34931_comb[31:8];
  assign p5_bit_slice_34978_comb = p5_sub_34932_comb[31:8];
  assign p5_bit_slice_34979_comb = p5_sub_34933_comb[31:8];
  assign p5_bit_slice_34980_comb = p5_sub_34934_comb[31:8];
  assign p5_sub_35005_comb = p5_add_34963_comb - {p5_add_34918_comb, p4_umul_34291[2:0]};
  assign p5_sub_35008_comb = {p5_add_34920_comb, p5_add_34826_comb[0]} - {p5_add_34922_comb, p5_add_34827_comb[2:0]};
  assign p5_sub_35027_comb = p5_add_35006_comb - {p5_add_34965_comb, p4_umul_34308[2:0]};
  assign p5_sub_35028_comb = {p5_add_34969_comb, p5_add_34888_comb[0]} - {p5_add_34971_comb, p5_add_34889_comb[2:0]};
  assign p5_bit_slice_35130_comb = p5_sub_35105_comb[31:8];
  assign p5_bit_slice_35131_comb = p5_sub_35106_comb[31:8];
  assign p5_bit_slice_35132_comb = p5_sub_35107_comb[31:8];
  assign p5_bit_slice_35133_comb = p5_sub_35108_comb[31:8];
  assign p5_bit_slice_35134_comb = p5_sub_35109_comb[31:8];
  assign p5_bit_slice_35135_comb = p5_sub_35110_comb[31:8];
  assign p5_bit_slice_35136_comb = p5_sub_35111_comb[31:8];
  assign p5_bit_slice_35137_comb = p5_sub_35112_comb[31:8];
  assign p5_sub_35280_comb = p5_add_35236_comb - p5_add_35237_comb;
  assign p5_sub_35281_comb = p5_add_35238_comb - p5_add_35239_comb;
  assign p5_sub_35282_comb = p5_add_35240_comb - p5_add_35241_comb;
  assign p5_sub_35283_comb = p5_add_35242_comb - p5_add_35243_comb;
  assign p5_bit_slice_35284_comb = p5_umul_35244_comb[31:2];
  assign p5_bit_slice_35285_comb = p5_umul_35245_comb[31:2];
  assign p5_bit_slice_35286_comb = p5_umul_35246_comb[31:2];
  assign p5_bit_slice_35287_comb = p5_umul_35247_comb[31:2];
  assign p5_sub_35352_comb = p5_add_35315_comb - p5_add_35316_comb;
  assign p5_sub_35354_comb = p5_add_35318_comb - p5_add_35319_comb;
  assign p5_sub_35356_comb = p5_add_35321_comb - p5_add_35322_comb;
  assign p5_sub_35358_comb = p5_add_35324_comb - p5_add_35325_comb;
  assign p5_add_35363_comb = p5_add_35288_comb[31:2] + {p5_add_35289_comb, p5_add_35138_comb[1:0], p4_umul_34389[4:2]};
  assign p5_sub_35366_comb = {p5_add_35294_comb, p4_umul_34273[2:0]} - {p5_add_35296_comb, p5_add_35208_comb[0], p4_umul_34306[0]};
  assign p5_sub_35369_comb = {p5_add_35303_comb, p4_umul_34306[0]} - {p5_add_35304_comb, p4_umul_34273[1:0]};
  assign p5_sub_35372_comb = {p5_add_35308_comb, p4_umul_34305[1:0]} - {p5_add_35310_comb, p4_umul_34273[1:0]};
  assign p5_bit_slice_35375_comb = p5_umul_35359_comb[31:5];
  assign p5_bit_slice_35376_comb = p5_umul_35360_comb[31:5];
  assign p5_bit_slice_35377_comb = p5_umul_35361_comb[31:5];
  assign p5_bit_slice_35378_comb = p5_umul_35362_comb[31:5];
  assign p5_add_35379_comb = p5_add_35332_comb[31:2] + {p5_add_35333_comb, p5_add_35178_comb[1:0], p4_umul_34412[4:2]};
  assign p5_sub_35380_comb = {p5_add_35337_comb, p4_umul_34285[2:0]} - {p5_add_35339_comb, p5_add_35260_comb[0], p4_umul_34316[0]};
  assign p5_sub_35381_comb = {p5_add_35344_comb, p4_umul_34316[0]} - {p5_add_35345_comb, p4_umul_34285[1:0]};
  assign p5_sub_35382_comb = {p5_add_35348_comb, p4_umul_34315[1:0]} - {p5_add_35350_comb, p4_umul_34285[1:0]};
  assign p5_add_35383_comb = p5_sign_ext_35180_comb + p5_sign_ext_35182_comb;
  assign p5_add_35384_comb = p5_sign_ext_35184_comb + p5_sign_ext_35186_comb;
  assign p5_add_35385_comb = p5_sign_ext_35188_comb + p5_sign_ext_35190_comb;
  assign p5_add_35386_comb = p5_sign_ext_35192_comb + p5_sign_ext_35194_comb;
  assign p5_add_35387_comb = p5_sign_ext_35181_comb + p5_sign_ext_35179_comb;
  assign p5_add_35388_comb = p5_sign_ext_35185_comb + p5_sign_ext_35183_comb;
  assign p5_add_35389_comb = p5_sign_ext_35189_comb + p5_sign_ext_35187_comb;
  assign p5_add_35390_comb = p5_sign_ext_35193_comb + p5_sign_ext_35191_comb;
  assign p5_umul_35351_comb = umul32b_32b_x_12b(p5_sign_ext_35157_comb, 12'hec8);
  assign p5_umul_35353_comb = umul32b_32b_x_12b(p5_sign_ext_35159_comb, 12'hec8);
  assign p5_umul_35355_comb = umul32b_32b_x_12b(p5_sign_ext_35161_comb, 12'hec8);
  assign p5_umul_35357_comb = umul32b_32b_x_12b(p5_sign_ext_35163_comb, 12'hec8);

  // Registers for pipe stage 5:
  reg [23:0] p5_bit_slice_34894;
  reg [23:0] p5_bit_slice_34895;
  reg [23:0] p5_bit_slice_34900;
  reg [23:0] p5_bit_slice_34901;
  reg [23:0] p5_bit_slice_34906;
  reg [23:0] p5_bit_slice_34907;
  reg [23:0] p5_bit_slice_34912;
  reg [23:0] p5_bit_slice_34913;
  reg [23:0] p5_bit_slice_34973;
  reg [23:0] p5_bit_slice_34974;
  reg [23:0] p5_bit_slice_34975;
  reg [23:0] p5_bit_slice_34976;
  reg [23:0] p5_bit_slice_34977;
  reg [23:0] p5_bit_slice_34978;
  reg [23:0] p5_bit_slice_34979;
  reg [23:0] p5_bit_slice_34980;
  reg [31:0] p5_sub_35005;
  reg [31:0] p5_sub_35008;
  reg [31:0] p5_sub_35027;
  reg [31:0] p5_sub_35028;
  reg [23:0] p5_bit_slice_35130;
  reg [23:0] p5_bit_slice_35131;
  reg [23:0] p5_bit_slice_35132;
  reg [23:0] p5_bit_slice_35133;
  reg [23:0] p5_bit_slice_35134;
  reg [23:0] p5_bit_slice_35135;
  reg [23:0] p5_bit_slice_35136;
  reg [23:0] p5_bit_slice_35137;
  reg [20:0] p5_bit_slice_33029;
  reg [20:0] p5_bit_slice_33030;
  reg [20:0] p5_bit_slice_33033;
  reg [20:0] p5_bit_slice_33034;
  reg [31:0] p5_sub_35280;
  reg [31:0] p5_sub_35281;
  reg [31:0] p5_sub_35282;
  reg [31:0] p5_sub_35283;
  reg [29:0] p5_bit_slice_35284;
  reg [29:0] p5_bit_slice_35285;
  reg [29:0] p5_bit_slice_35286;
  reg [29:0] p5_bit_slice_35287;
  reg [31:0] p5_sub_35352;
  reg [31:0] p5_sub_35354;
  reg [31:0] p5_sub_35356;
  reg [31:0] p5_sub_35358;
  reg [29:0] p5_add_35363;
  reg [31:0] p5_sub_35366;
  reg [31:0] p5_sub_35369;
  reg [31:0] p5_sub_35372;
  reg [26:0] p5_bit_slice_35375;
  reg [26:0] p5_bit_slice_35376;
  reg [26:0] p5_bit_slice_35377;
  reg [26:0] p5_bit_slice_35378;
  reg [29:0] p5_add_35379;
  reg [31:0] p5_sub_35380;
  reg [31:0] p5_sub_35381;
  reg [31:0] p5_sub_35382;
  reg [31:0] p5_add_35383;
  reg [31:0] p5_add_35384;
  reg [31:0] p5_add_35385;
  reg [31:0] p5_add_35386;
  reg [31:0] p5_add_35387;
  reg [31:0] p5_add_35388;
  reg [31:0] p5_add_35389;
  reg [31:0] p5_add_35390;
  reg [31:0] p5_umul_34389;
  reg [31:0] p5_umul_34412;
  reg [31:0] p5_umul_34413;
  reg [31:0] p5_umul_34416;
  reg [31:0] p5_umul_35351;
  reg [31:0] p5_umul_35353;
  reg [31:0] p5_umul_35355;
  reg [31:0] p5_umul_35357;
  always_ff @ (posedge clk) begin
    p5_bit_slice_34894 <= p5_bit_slice_34894_comb;
    p5_bit_slice_34895 <= p5_bit_slice_34895_comb;
    p5_bit_slice_34900 <= p5_bit_slice_34900_comb;
    p5_bit_slice_34901 <= p5_bit_slice_34901_comb;
    p5_bit_slice_34906 <= p5_bit_slice_34906_comb;
    p5_bit_slice_34907 <= p5_bit_slice_34907_comb;
    p5_bit_slice_34912 <= p5_bit_slice_34912_comb;
    p5_bit_slice_34913 <= p5_bit_slice_34913_comb;
    p5_bit_slice_34973 <= p5_bit_slice_34973_comb;
    p5_bit_slice_34974 <= p5_bit_slice_34974_comb;
    p5_bit_slice_34975 <= p5_bit_slice_34975_comb;
    p5_bit_slice_34976 <= p5_bit_slice_34976_comb;
    p5_bit_slice_34977 <= p5_bit_slice_34977_comb;
    p5_bit_slice_34978 <= p5_bit_slice_34978_comb;
    p5_bit_slice_34979 <= p5_bit_slice_34979_comb;
    p5_bit_slice_34980 <= p5_bit_slice_34980_comb;
    p5_sub_35005 <= p5_sub_35005_comb;
    p5_sub_35008 <= p5_sub_35008_comb;
    p5_sub_35027 <= p5_sub_35027_comb;
    p5_sub_35028 <= p5_sub_35028_comb;
    p5_bit_slice_35130 <= p5_bit_slice_35130_comb;
    p5_bit_slice_35131 <= p5_bit_slice_35131_comb;
    p5_bit_slice_35132 <= p5_bit_slice_35132_comb;
    p5_bit_slice_35133 <= p5_bit_slice_35133_comb;
    p5_bit_slice_35134 <= p5_bit_slice_35134_comb;
    p5_bit_slice_35135 <= p5_bit_slice_35135_comb;
    p5_bit_slice_35136 <= p5_bit_slice_35136_comb;
    p5_bit_slice_35137 <= p5_bit_slice_35137_comb;
    p5_bit_slice_33029 <= p4_bit_slice_33029;
    p5_bit_slice_33030 <= p4_bit_slice_33030;
    p5_bit_slice_33033 <= p4_bit_slice_33033;
    p5_bit_slice_33034 <= p4_bit_slice_33034;
    p5_sub_35280 <= p5_sub_35280_comb;
    p5_sub_35281 <= p5_sub_35281_comb;
    p5_sub_35282 <= p5_sub_35282_comb;
    p5_sub_35283 <= p5_sub_35283_comb;
    p5_bit_slice_35284 <= p5_bit_slice_35284_comb;
    p5_bit_slice_35285 <= p5_bit_slice_35285_comb;
    p5_bit_slice_35286 <= p5_bit_slice_35286_comb;
    p5_bit_slice_35287 <= p5_bit_slice_35287_comb;
    p5_sub_35352 <= p5_sub_35352_comb;
    p5_sub_35354 <= p5_sub_35354_comb;
    p5_sub_35356 <= p5_sub_35356_comb;
    p5_sub_35358 <= p5_sub_35358_comb;
    p5_add_35363 <= p5_add_35363_comb;
    p5_sub_35366 <= p5_sub_35366_comb;
    p5_sub_35369 <= p5_sub_35369_comb;
    p5_sub_35372 <= p5_sub_35372_comb;
    p5_bit_slice_35375 <= p5_bit_slice_35375_comb;
    p5_bit_slice_35376 <= p5_bit_slice_35376_comb;
    p5_bit_slice_35377 <= p5_bit_slice_35377_comb;
    p5_bit_slice_35378 <= p5_bit_slice_35378_comb;
    p5_add_35379 <= p5_add_35379_comb;
    p5_sub_35380 <= p5_sub_35380_comb;
    p5_sub_35381 <= p5_sub_35381_comb;
    p5_sub_35382 <= p5_sub_35382_comb;
    p5_add_35383 <= p5_add_35383_comb;
    p5_add_35384 <= p5_add_35384_comb;
    p5_add_35385 <= p5_add_35385_comb;
    p5_add_35386 <= p5_add_35386_comb;
    p5_add_35387 <= p5_add_35387_comb;
    p5_add_35388 <= p5_add_35388_comb;
    p5_add_35389 <= p5_add_35389_comb;
    p5_add_35390 <= p5_add_35390_comb;
    p5_umul_34389 <= p4_umul_34389;
    p5_umul_34412 <= p4_umul_34412;
    p5_umul_34413 <= p4_umul_34413;
    p5_umul_34416 <= p4_umul_34416;
    p5_umul_35351 <= p5_umul_35351_comb;
    p5_umul_35353 <= p5_umul_35353_comb;
    p5_umul_35355 <= p5_umul_35355_comb;
    p5_umul_35357 <= p5_umul_35357_comb;
  end

  // ===== Pipe stage 6:
  wire [29:0] p6_add_35651_comb;
  wire [29:0] p6_add_35653_comb;
  wire [29:0] p6_add_35655_comb;
  wire [29:0] p6_add_35657_comb;
  wire [26:0] p6_add_35707_comb;
  wire [26:0] p6_add_35709_comb;
  wire [26:0] p6_add_35711_comb;
  wire [26:0] p6_add_35713_comb;
  wire [28:0] p6_concat_35731_comb;
  wire [18:0] p6_add_35715_comb;
  wire [4:0] p6_bit_slice_35716_comb;
  wire [28:0] p6_concat_35732_comb;
  wire [18:0] p6_add_35718_comb;
  wire [4:0] p6_bit_slice_35719_comb;
  wire [28:0] p6_concat_35733_comb;
  wire [18:0] p6_add_35721_comb;
  wire [4:0] p6_bit_slice_35722_comb;
  wire [28:0] p6_concat_35734_comb;
  wire [18:0] p6_add_35724_comb;
  wire [4:0] p6_bit_slice_35725_comb;
  wire [31:0] p6_sign_ext_35743_comb;
  wire [23:0] p6_bit_slice_35717_comb;
  wire [31:0] p6_sign_ext_35745_comb;
  wire [23:0] p6_bit_slice_35720_comb;
  wire [31:0] p6_sign_ext_35747_comb;
  wire [23:0] p6_bit_slice_35723_comb;
  wire [31:0] p6_sign_ext_35749_comb;
  wire [23:0] p6_bit_slice_35726_comb;
  wire [18:0] p6_add_35751_comb;
  wire [18:0] p6_add_35753_comb;
  wire [18:0] p6_add_35755_comb;
  wire [18:0] p6_add_35757_comb;
  wire [23:0] p6_add_35760_comb;
  wire [23:0] p6_add_35762_comb;
  wire [23:0] p6_add_35764_comb;
  wire [23:0] p6_add_35766_comb;
  wire [23:0] p6_bit_slice_35767_comb;
  wire [23:0] p6_bit_slice_35768_comb;
  wire [23:0] p6_bit_slice_35769_comb;
  wire [23:0] p6_bit_slice_35770_comb;
  wire [31:0] p6_sign_ext_35535_comb;
  wire [31:0] p6_sign_ext_35536_comb;
  wire [31:0] p6_sign_ext_35537_comb;
  wire [31:0] p6_sign_ext_35538_comb;
  wire [31:0] p6_sign_ext_35539_comb;
  wire [31:0] p6_sign_ext_35540_comb;
  wire [31:0] p6_sign_ext_35541_comb;
  wire [31:0] p6_sign_ext_35542_comb;
  wire [23:0] p6_add_35779_comb;
  wire [23:0] p6_add_35781_comb;
  wire [23:0] p6_add_35783_comb;
  wire [23:0] p6_add_35785_comb;
  wire [23:0] p6_add_35791_comb;
  wire [23:0] p6_add_35793_comb;
  wire [23:0] p6_add_35795_comb;
  wire [23:0] p6_add_35797_comb;
  wire [31:0] p6_add_35543_comb;
  wire [31:0] p6_add_35545_comb;
  wire [31:0] p6_add_35547_comb;
  wire [31:0] p6_add_35549_comb;
  wire [31:0] p6_concat_35799_comb;
  wire [31:0] p6_concat_35800_comb;
  wire [31:0] p6_concat_35801_comb;
  wire [31:0] p6_concat_35802_comb;
  wire [31:0] p6_sub_35803_comb;
  wire [31:0] p6_sub_35804_comb;
  wire [31:0] p6_sub_35805_comb;
  wire [31:0] p6_sub_35806_comb;
  wire [31:0] p6_add_35808_comb;
  wire [31:0] p6_add_35810_comb;
  wire [31:0] p6_add_35812_comb;
  wire [31:0] p6_add_35814_comb;
  wire [31:0] p6_umul_35565_comb;
  wire [31:0] p6_umul_35567_comb;
  wire [31:0] p6_umul_35587_comb;
  wire [31:0] p6_umul_35590_comb;
  wire [31:0] p6_umul_35647_comb;
  wire [31:0] p6_umul_35648_comb;
  wire [31:0] p6_umul_35649_comb;
  wire [31:0] p6_umul_35650_comb;
  wire [31:0] p6_umul_35680_comb;
  wire [31:0] p6_umul_35682_comb;
  wire [31:0] p6_umul_35684_comb;
  wire [31:0] p6_umul_35686_comb;
  wire [31:0] p6_sign_ext_35553_comb;
  wire [31:0] p6_sign_ext_35554_comb;
  wire [31:0] p6_sign_ext_35556_comb;
  wire [31:0] p6_sign_ext_35557_comb;
  wire [31:0] p6_sign_ext_35559_comb;
  wire [31:0] p6_sign_ext_35560_comb;
  wire [31:0] p6_sign_ext_35562_comb;
  wire [31:0] p6_sign_ext_35563_comb;
  wire [31:0] p6_umul_35555_comb;
  wire [31:0] p6_umul_35558_comb;
  wire [31:0] p6_umul_35561_comb;
  wire [31:0] p6_umul_35564_comb;
  wire [31:0] p6_umul_35591_comb;
  wire [31:0] p6_umul_35597_comb;
  wire [31:0] p6_umul_35603_comb;
  wire [31:0] p6_umul_35609_comb;
  wire [31:0] p6_add_35815_comb;
  wire [31:0] p6_add_35816_comb;
  wire [31:0] p6_add_35817_comb;
  wire [31:0] p6_add_35818_comb;
  wire [31:0] p6_add_35819_comb;
  wire [31:0] p6_add_35820_comb;
  wire [31:0] p6_add_35821_comb;
  wire [31:0] p6_add_35822_comb;
  wire [31:0] p6_sub_35823_comb;
  wire [31:0] p6_sub_35824_comb;
  wire [31:0] p6_sub_35825_comb;
  wire [31:0] p6_sub_35826_comb;
  wire [31:0] p6_sub_35827_comb;
  wire [31:0] p6_sub_35828_comb;
  wire [31:0] p6_sub_35829_comb;
  wire [31:0] p6_sub_35830_comb;
  wire [31:0] p6_add_35570_comb;
  wire [31:0] p6_add_35574_comb;
  wire [31:0] p6_add_35578_comb;
  wire [31:0] p6_add_35582_comb;
  wire [29:0] p6_bit_slice_35572_comb;
  wire [29:0] p6_bit_slice_35576_comb;
  wire [29:0] p6_bit_slice_35580_comb;
  wire [29:0] p6_bit_slice_35584_comb;
  wire [1:0] p6_bit_slice_35595_comb;
  wire [1:0] p6_bit_slice_35601_comb;
  wire [1:0] p6_bit_slice_35607_comb;
  wire [1:0] p6_bit_slice_35613_comb;
  wire [29:0] p6_bit_slice_35621_comb;
  wire [29:0] p6_bit_slice_35625_comb;
  wire [29:0] p6_bit_slice_35629_comb;
  wire [29:0] p6_bit_slice_35633_comb;
  wire [31:0] p6_sub_35679_comb;
  wire [31:0] p6_sub_35681_comb;
  wire [31:0] p6_sub_35683_comb;
  wire [31:0] p6_sub_35685_comb;
  wire [17:0] p6_bit_slice_35831_comb;
  wire [17:0] p6_bit_slice_35832_comb;
  wire [17:0] p6_bit_slice_35833_comb;
  wire [17:0] p6_bit_slice_35834_comb;
  wire [17:0] p6_bit_slice_35835_comb;
  wire [17:0] p6_bit_slice_35836_comb;
  wire [17:0] p6_bit_slice_35837_comb;
  wire [17:0] p6_bit_slice_35838_comb;
  wire [17:0] p6_bit_slice_35839_comb;
  wire [17:0] p6_bit_slice_35840_comb;
  wire [17:0] p6_bit_slice_35841_comb;
  wire [17:0] p6_bit_slice_35842_comb;
  wire [17:0] p6_bit_slice_35843_comb;
  wire [17:0] p6_bit_slice_35844_comb;
  wire [17:0] p6_bit_slice_35845_comb;
  wire [17:0] p6_bit_slice_35846_comb;
  wire [24:0] p6_add_35615_comb;
  wire [24:0] p6_add_35618_comb;
  wire [24:0] p6_add_35637_comb;
  wire [24:0] p6_add_35638_comb;
  wire [24:0] p6_add_35675_comb;
  wire [24:0] p6_add_35676_comb;
  wire [24:0] p6_add_35677_comb;
  wire [24:0] p6_add_35678_comb;
  wire [24:0] p6_add_35727_comb;
  wire [24:0] p6_add_35728_comb;
  wire [24:0] p6_add_35729_comb;
  wire [24:0] p6_add_35730_comb;
  wire [31:0] p6_umul_35592_comb;
  wire [31:0] p6_umul_35598_comb;
  wire [31:0] p6_umul_35604_comb;
  wire [31:0] p6_umul_35610_comb;
  wire [31:0] p6_umul_35622_comb;
  wire [31:0] p6_umul_35623_comb;
  wire [31:0] p6_umul_35624_comb;
  wire [31:0] p6_umul_35626_comb;
  wire [31:0] p6_umul_35627_comb;
  wire [31:0] p6_umul_35628_comb;
  wire [31:0] p6_umul_35630_comb;
  wire [31:0] p6_umul_35631_comb;
  wire [31:0] p6_umul_35632_comb;
  wire [31:0] p6_umul_35634_comb;
  wire [31:0] p6_umul_35635_comb;
  wire [31:0] p6_umul_35636_comb;
  assign p6_add_35651_comb = p5_bit_slice_35284 + 30'h0000_0001;
  assign p6_add_35653_comb = p5_bit_slice_35285 + 30'h0000_0001;
  assign p6_add_35655_comb = p5_bit_slice_35286 + 30'h0000_0001;
  assign p6_add_35657_comb = p5_bit_slice_35287 + 30'h0000_0001;
  assign p6_add_35707_comb = p5_bit_slice_35375 + p6_add_35651_comb[29:3];
  assign p6_add_35709_comb = p5_bit_slice_35376 + p6_add_35653_comb[29:3];
  assign p6_add_35711_comb = p5_bit_slice_35377 + p6_add_35655_comb[29:3];
  assign p6_add_35713_comb = p5_bit_slice_35378 + p6_add_35657_comb[29:3];
  assign p6_concat_35731_comb = {p6_add_35707_comb, p6_add_35651_comb[2:1]};
  assign p6_add_35715_comb = p5_add_35363[29:11] + 19'h0_0001;
  assign p6_bit_slice_35716_comb = p5_add_35363[10:6];
  assign p6_concat_35732_comb = {p6_add_35709_comb, p6_add_35653_comb[2:1]};
  assign p6_add_35718_comb = p5_sub_35366[31:13] + 19'h0_0001;
  assign p6_bit_slice_35719_comb = p5_sub_35366[12:8];
  assign p6_concat_35733_comb = {p6_add_35711_comb, p6_add_35655_comb[2:1]};
  assign p6_add_35721_comb = p5_sub_35369[31:13] + 19'h0_0001;
  assign p6_bit_slice_35722_comb = p5_sub_35369[12:8];
  assign p6_concat_35734_comb = {p6_add_35713_comb, p6_add_35657_comb[2:1]};
  assign p6_add_35724_comb = p5_sub_35372[31:13] + 19'h0_0001;
  assign p6_bit_slice_35725_comb = p5_sub_35372[12:8];
  assign p6_sign_ext_35743_comb = {{3{p6_concat_35731_comb[28]}}, p6_concat_35731_comb};
  assign p6_bit_slice_35717_comb = p5_add_35379[29:6];
  assign p6_sign_ext_35745_comb = {{3{p6_concat_35732_comb[28]}}, p6_concat_35732_comb};
  assign p6_bit_slice_35720_comb = p5_sub_35380[31:8];
  assign p6_sign_ext_35747_comb = {{3{p6_concat_35733_comb[28]}}, p6_concat_35733_comb};
  assign p6_bit_slice_35723_comb = p5_sub_35381[31:8];
  assign p6_sign_ext_35749_comb = {{3{p6_concat_35734_comb[28]}}, p6_concat_35734_comb};
  assign p6_bit_slice_35726_comb = p5_sub_35382[31:8];
  assign p6_add_35751_comb = p5_add_35379[29:11] + 19'h0_0001;
  assign p6_add_35753_comb = p5_sub_35380[31:13] + 19'h0_0001;
  assign p6_add_35755_comb = p5_sub_35381[31:13] + 19'h0_0001;
  assign p6_add_35757_comb = p5_sub_35382[31:13] + 19'h0_0001;
  assign p6_add_35760_comb = p6_bit_slice_35717_comb + {p6_add_35715_comb, p6_bit_slice_35716_comb};
  assign p6_add_35762_comb = p6_bit_slice_35720_comb + {p6_add_35718_comb, p6_bit_slice_35719_comb};
  assign p6_add_35764_comb = p6_bit_slice_35723_comb + {p6_add_35721_comb, p6_bit_slice_35722_comb};
  assign p6_add_35766_comb = p6_bit_slice_35726_comb + {p6_add_35724_comb, p6_bit_slice_35725_comb};
  assign p6_bit_slice_35767_comb = p5_add_35363[29:6];
  assign p6_bit_slice_35768_comb = p5_sub_35366[31:8];
  assign p6_bit_slice_35769_comb = p5_sub_35369[31:8];
  assign p6_bit_slice_35770_comb = p5_sub_35372[31:8];
  assign p6_sign_ext_35535_comb = {{8{p5_bit_slice_34894[23]}}, p5_bit_slice_34894};
  assign p6_sign_ext_35536_comb = {{8{p5_bit_slice_34895[23]}}, p5_bit_slice_34895};
  assign p6_sign_ext_35537_comb = {{8{p5_bit_slice_34900[23]}}, p5_bit_slice_34900};
  assign p6_sign_ext_35538_comb = {{8{p5_bit_slice_34901[23]}}, p5_bit_slice_34901};
  assign p6_sign_ext_35539_comb = {{8{p5_bit_slice_34906[23]}}, p5_bit_slice_34906};
  assign p6_sign_ext_35540_comb = {{8{p5_bit_slice_34907[23]}}, p5_bit_slice_34907};
  assign p6_sign_ext_35541_comb = {{8{p5_bit_slice_34912[23]}}, p5_bit_slice_34912};
  assign p6_sign_ext_35542_comb = {{8{p5_bit_slice_34913[23]}}, p5_bit_slice_34913};
  assign p6_add_35779_comb = p6_sign_ext_35743_comb[31:8] + p6_add_35760_comb;
  assign p6_add_35781_comb = p6_sign_ext_35745_comb[31:8] + p6_add_35762_comb;
  assign p6_add_35783_comb = p6_sign_ext_35747_comb[31:8] + p6_add_35764_comb;
  assign p6_add_35785_comb = p6_sign_ext_35749_comb[31:8] + p6_add_35766_comb;
  assign p6_add_35791_comb = {p6_add_35751_comb, p5_add_35379[10:6]} + p6_bit_slice_35767_comb;
  assign p6_add_35793_comb = {p6_add_35753_comb, p5_sub_35380[12:8]} + p6_bit_slice_35768_comb;
  assign p6_add_35795_comb = {p6_add_35755_comb, p5_sub_35381[12:8]} + p6_bit_slice_35769_comb;
  assign p6_add_35797_comb = {p6_add_35757_comb, p5_sub_35382[12:8]} + p6_bit_slice_35770_comb;
  assign p6_add_35543_comb = p6_sign_ext_35535_comb + p6_sign_ext_35536_comb;
  assign p6_add_35545_comb = p6_sign_ext_35537_comb + p6_sign_ext_35538_comb;
  assign p6_add_35547_comb = p6_sign_ext_35539_comb + p6_sign_ext_35540_comb;
  assign p6_add_35549_comb = p6_sign_ext_35541_comb + p6_sign_ext_35542_comb;
  assign p6_concat_35799_comb = {p6_add_35779_comb, p6_add_35707_comb[5:0], p6_add_35651_comb[2:1]};
  assign p6_concat_35800_comb = {p6_add_35781_comb, p6_add_35709_comb[5:0], p6_add_35653_comb[2:1]};
  assign p6_concat_35801_comb = {p6_add_35783_comb, p6_add_35711_comb[5:0], p6_add_35655_comb[2:1]};
  assign p6_concat_35802_comb = {p6_add_35785_comb, p6_add_35713_comb[5:0], p6_add_35657_comb[2:1]};
  assign p6_sub_35803_comb = {p6_add_35760_comb, 8'h00} - p6_sign_ext_35743_comb;
  assign p6_sub_35804_comb = {p6_add_35762_comb, 8'h00} - p6_sign_ext_35745_comb;
  assign p6_sub_35805_comb = {p6_add_35764_comb, 8'h00} - p6_sign_ext_35747_comb;
  assign p6_sub_35806_comb = {p6_add_35766_comb, 8'h00} - p6_sign_ext_35749_comb;
  assign p6_add_35808_comb = p6_sign_ext_35743_comb + p5_add_35383;
  assign p6_add_35810_comb = p6_sign_ext_35745_comb + p5_add_35384;
  assign p6_add_35812_comb = p6_sign_ext_35747_comb + p5_add_35385;
  assign p6_add_35814_comb = p6_sign_ext_35749_comb + p5_add_35386;
  assign p6_umul_35565_comb = umul32b_32b_x_8b(p5_sub_35005, 8'hb5);
  assign p6_umul_35567_comb = umul32b_32b_x_8b(p5_sub_35008, 8'hb5);
  assign p6_umul_35587_comb = umul32b_32b_x_8b(p5_sub_35027, 8'hb5);
  assign p6_umul_35590_comb = umul32b_32b_x_8b(p5_sub_35028, 8'hb5);
  assign p6_umul_35647_comb = umul32b_32b_x_8b(p5_sub_35280, 8'hb5);
  assign p6_umul_35648_comb = umul32b_32b_x_8b(p5_sub_35281, 8'hb5);
  assign p6_umul_35649_comb = umul32b_32b_x_8b(p5_sub_35282, 8'hb5);
  assign p6_umul_35650_comb = umul32b_32b_x_8b(p5_sub_35283, 8'hb5);
  assign p6_umul_35680_comb = umul32b_32b_x_8b(p5_sub_35352, 8'hb5);
  assign p6_umul_35682_comb = umul32b_32b_x_8b(p5_sub_35354, 8'hb5);
  assign p6_umul_35684_comb = umul32b_32b_x_8b(p5_sub_35356, 8'hb5);
  assign p6_umul_35686_comb = umul32b_32b_x_8b(p5_sub_35358, 8'hb5);
  assign p6_sign_ext_35553_comb = {{8{p5_bit_slice_34973[23]}}, p5_bit_slice_34973};
  assign p6_sign_ext_35554_comb = {{8{p5_bit_slice_34974[23]}}, p5_bit_slice_34974};
  assign p6_sign_ext_35556_comb = {{8{p5_bit_slice_34975[23]}}, p5_bit_slice_34975};
  assign p6_sign_ext_35557_comb = {{8{p5_bit_slice_34976[23]}}, p5_bit_slice_34976};
  assign p6_sign_ext_35559_comb = {{8{p5_bit_slice_34977[23]}}, p5_bit_slice_34977};
  assign p6_sign_ext_35560_comb = {{8{p5_bit_slice_34978[23]}}, p5_bit_slice_34978};
  assign p6_sign_ext_35562_comb = {{8{p5_bit_slice_34979[23]}}, p5_bit_slice_34979};
  assign p6_sign_ext_35563_comb = {{8{p5_bit_slice_34980[23]}}, p5_bit_slice_34980};
  assign p6_umul_35555_comb = umul32b_32b_x_10b(p6_add_35543_comb, 10'h235);
  assign p6_umul_35558_comb = umul32b_32b_x_10b(p6_add_35545_comb, 10'h235);
  assign p6_umul_35561_comb = umul32b_32b_x_10b(p6_add_35547_comb, 10'h235);
  assign p6_umul_35564_comb = umul32b_32b_x_10b(p6_add_35549_comb, 10'h235);
  assign p6_umul_35591_comb = umul32b_32b_x_12b(p6_sign_ext_35535_comb, 12'h8e4);
  assign p6_umul_35597_comb = umul32b_32b_x_12b(p6_sign_ext_35537_comb, 12'h8e4);
  assign p6_umul_35603_comb = umul32b_32b_x_12b(p6_sign_ext_35539_comb, 12'h8e4);
  assign p6_umul_35609_comb = umul32b_32b_x_12b(p6_sign_ext_35541_comb, 12'h8e4);
  assign p6_add_35815_comb = p5_add_35387 + p6_concat_35799_comb;
  assign p6_add_35816_comb = p5_add_35388 + p6_concat_35800_comb;
  assign p6_add_35817_comb = p5_add_35389 + p6_concat_35801_comb;
  assign p6_add_35818_comb = p5_add_35390 + p6_concat_35802_comb;
  assign p6_add_35819_comb = p6_sub_35803_comb + p5_add_35383;
  assign p6_add_35820_comb = p6_sub_35804_comb + p5_add_35384;
  assign p6_add_35821_comb = p6_sub_35805_comb + p5_add_35385;
  assign p6_add_35822_comb = p6_sub_35806_comb + p5_add_35386;
  assign p6_sub_35823_comb = {p6_add_35791_comb, 8'h00} - p6_add_35808_comb;
  assign p6_sub_35824_comb = {p6_add_35793_comb, 8'h00} - p6_add_35810_comb;
  assign p6_sub_35825_comb = {p6_add_35795_comb, 8'h00} - p6_add_35812_comb;
  assign p6_sub_35826_comb = {p6_add_35797_comb, 8'h00} - p6_add_35814_comb;
  assign p6_sub_35827_comb = p6_concat_35799_comb - p5_add_35387;
  assign p6_sub_35828_comb = p6_concat_35800_comb - p5_add_35388;
  assign p6_sub_35829_comb = p6_concat_35801_comb - p5_add_35389;
  assign p6_sub_35830_comb = p6_concat_35802_comb - p5_add_35390;
  assign p6_add_35570_comb = p6_sign_ext_35553_comb + p6_sign_ext_35554_comb;
  assign p6_add_35574_comb = p6_sign_ext_35556_comb + p6_sign_ext_35557_comb;
  assign p6_add_35578_comb = p6_sign_ext_35559_comb + p6_sign_ext_35560_comb;
  assign p6_add_35582_comb = p6_sign_ext_35562_comb + p6_sign_ext_35563_comb;
  assign p6_bit_slice_35572_comb = p6_umul_35555_comb[31:2];
  assign p6_bit_slice_35576_comb = p6_umul_35558_comb[31:2];
  assign p6_bit_slice_35580_comb = p6_umul_35561_comb[31:2];
  assign p6_bit_slice_35584_comb = p6_umul_35564_comb[31:2];
  assign p6_bit_slice_35595_comb = p6_umul_35555_comb[1:0];
  assign p6_bit_slice_35601_comb = p6_umul_35558_comb[1:0];
  assign p6_bit_slice_35607_comb = p6_umul_35561_comb[1:0];
  assign p6_bit_slice_35613_comb = p6_umul_35564_comb[1:0];
  assign p6_bit_slice_35621_comb = p6_umul_35591_comb[31:2];
  assign p6_bit_slice_35625_comb = p6_umul_35597_comb[31:2];
  assign p6_bit_slice_35629_comb = p6_umul_35603_comb[31:2];
  assign p6_bit_slice_35633_comb = p6_umul_35609_comb[31:2];
  assign p6_sub_35679_comb = {p6_add_35651_comb, 2'h0} - p5_umul_35351;
  assign p6_sub_35681_comb = {p6_add_35653_comb, 2'h0} - p5_umul_35353;
  assign p6_sub_35683_comb = {p6_add_35655_comb, 2'h0} - p5_umul_35355;
  assign p6_sub_35685_comb = {p6_add_35657_comb, 2'h0} - p5_umul_35357;
  assign p6_bit_slice_35831_comb = p6_add_35815_comb[31:14];
  assign p6_bit_slice_35832_comb = p6_add_35816_comb[31:14];
  assign p6_bit_slice_35833_comb = p6_add_35817_comb[31:14];
  assign p6_bit_slice_35834_comb = p6_add_35818_comb[31:14];
  assign p6_bit_slice_35835_comb = p6_add_35819_comb[31:14];
  assign p6_bit_slice_35836_comb = p6_add_35820_comb[31:14];
  assign p6_bit_slice_35837_comb = p6_add_35821_comb[31:14];
  assign p6_bit_slice_35838_comb = p6_add_35822_comb[31:14];
  assign p6_bit_slice_35839_comb = p6_sub_35823_comb[31:14];
  assign p6_bit_slice_35840_comb = p6_sub_35824_comb[31:14];
  assign p6_bit_slice_35841_comb = p6_sub_35825_comb[31:14];
  assign p6_bit_slice_35842_comb = p6_sub_35826_comb[31:14];
  assign p6_bit_slice_35843_comb = p6_sub_35827_comb[31:14];
  assign p6_bit_slice_35844_comb = p6_sub_35828_comb[31:14];
  assign p6_bit_slice_35845_comb = p6_sub_35829_comb[31:14];
  assign p6_bit_slice_35846_comb = p6_sub_35830_comb[31:14];
  assign p6_add_35615_comb = p6_umul_35565_comb[31:7] + 25'h000_0001;
  assign p6_add_35618_comb = p6_umul_35567_comb[31:7] + 25'h000_0001;
  assign p6_add_35637_comb = p6_umul_35587_comb[31:7] + 25'h000_0001;
  assign p6_add_35638_comb = p6_umul_35590_comb[31:7] + 25'h000_0001;
  assign p6_add_35675_comb = p6_umul_35647_comb[31:7] + 25'h000_0001;
  assign p6_add_35676_comb = p6_umul_35648_comb[31:7] + 25'h000_0001;
  assign p6_add_35677_comb = p6_umul_35649_comb[31:7] + 25'h000_0001;
  assign p6_add_35678_comb = p6_umul_35650_comb[31:7] + 25'h000_0001;
  assign p6_add_35727_comb = p6_umul_35680_comb[31:7] + 25'h000_0001;
  assign p6_add_35728_comb = p6_umul_35682_comb[31:7] + 25'h000_0001;
  assign p6_add_35729_comb = p6_umul_35684_comb[31:7] + 25'h000_0001;
  assign p6_add_35730_comb = p6_umul_35686_comb[31:7] + 25'h000_0001;
  assign p6_umul_35592_comb = umul32b_32b_x_12b(p6_add_35570_comb, 12'h968);
  assign p6_umul_35598_comb = umul32b_32b_x_12b(p6_add_35574_comb, 12'h968);
  assign p6_umul_35604_comb = umul32b_32b_x_12b(p6_add_35578_comb, 12'h968);
  assign p6_umul_35610_comb = umul32b_32b_x_12b(p6_add_35582_comb, 12'h968);
  assign p6_umul_35622_comb = umul32b_32b_x_12b(p6_sign_ext_35554_comb, 12'hfb1);
  assign p6_umul_35623_comb = umul32b_32b_x_10b(p6_sign_ext_35553_comb, 10'h31f);
  assign p6_umul_35624_comb = umul32b_32b_x_12b(p6_sign_ext_35536_comb, 12'hd4e);
  assign p6_umul_35626_comb = umul32b_32b_x_12b(p6_sign_ext_35557_comb, 12'hfb1);
  assign p6_umul_35627_comb = umul32b_32b_x_10b(p6_sign_ext_35556_comb, 10'h31f);
  assign p6_umul_35628_comb = umul32b_32b_x_12b(p6_sign_ext_35538_comb, 12'hd4e);
  assign p6_umul_35630_comb = umul32b_32b_x_12b(p6_sign_ext_35560_comb, 12'hfb1);
  assign p6_umul_35631_comb = umul32b_32b_x_10b(p6_sign_ext_35559_comb, 10'h31f);
  assign p6_umul_35632_comb = umul32b_32b_x_12b(p6_sign_ext_35540_comb, 12'hd4e);
  assign p6_umul_35634_comb = umul32b_32b_x_12b(p6_sign_ext_35563_comb, 12'hfb1);
  assign p6_umul_35635_comb = umul32b_32b_x_10b(p6_sign_ext_35562_comb, 10'h31f);
  assign p6_umul_35636_comb = umul32b_32b_x_12b(p6_sign_ext_35542_comb, 12'hd4e);

  // Registers for pipe stage 6:
  reg [29:0] p6_bit_slice_35572;
  reg [29:0] p6_bit_slice_35576;
  reg [29:0] p6_bit_slice_35580;
  reg [29:0] p6_bit_slice_35584;
  reg [1:0] p6_bit_slice_35595;
  reg [1:0] p6_bit_slice_35601;
  reg [1:0] p6_bit_slice_35607;
  reg [1:0] p6_bit_slice_35613;
  reg [29:0] p6_bit_slice_35621;
  reg [29:0] p6_bit_slice_35625;
  reg [29:0] p6_bit_slice_35629;
  reg [29:0] p6_bit_slice_35633;
  reg [23:0] p6_bit_slice_35130;
  reg [23:0] p6_bit_slice_35131;
  reg [23:0] p6_bit_slice_35132;
  reg [23:0] p6_bit_slice_35133;
  reg [23:0] p6_bit_slice_35134;
  reg [23:0] p6_bit_slice_35135;
  reg [23:0] p6_bit_slice_35136;
  reg [23:0] p6_bit_slice_35137;
  reg [20:0] p6_bit_slice_33029;
  reg [20:0] p6_bit_slice_33030;
  reg [20:0] p6_bit_slice_33033;
  reg [20:0] p6_bit_slice_33034;
  reg [31:0] p6_sub_35679;
  reg [31:0] p6_sub_35681;
  reg [31:0] p6_sub_35683;
  reg [31:0] p6_sub_35685;
  reg [4:0] p6_bit_slice_35716;
  reg [23:0] p6_bit_slice_35717;
  reg [4:0] p6_bit_slice_35719;
  reg [23:0] p6_bit_slice_35720;
  reg [4:0] p6_bit_slice_35722;
  reg [23:0] p6_bit_slice_35723;
  reg [4:0] p6_bit_slice_35725;
  reg [23:0] p6_bit_slice_35726;
  reg [23:0] p6_bit_slice_35767;
  reg [23:0] p6_bit_slice_35768;
  reg [23:0] p6_bit_slice_35769;
  reg [23:0] p6_bit_slice_35770;
  reg [17:0] p6_bit_slice_35831;
  reg [17:0] p6_bit_slice_35832;
  reg [17:0] p6_bit_slice_35833;
  reg [17:0] p6_bit_slice_35834;
  reg [17:0] p6_bit_slice_35835;
  reg [17:0] p6_bit_slice_35836;
  reg [17:0] p6_bit_slice_35837;
  reg [17:0] p6_bit_slice_35838;
  reg [17:0] p6_bit_slice_35839;
  reg [17:0] p6_bit_slice_35840;
  reg [17:0] p6_bit_slice_35841;
  reg [17:0] p6_bit_slice_35842;
  reg [17:0] p6_bit_slice_35843;
  reg [17:0] p6_bit_slice_35844;
  reg [17:0] p6_bit_slice_35845;
  reg [17:0] p6_bit_slice_35846;
  reg [24:0] p6_add_35615;
  reg [24:0] p6_add_35618;
  reg [24:0] p6_add_35637;
  reg [24:0] p6_add_35638;
  reg [24:0] p6_add_35675;
  reg [24:0] p6_add_35676;
  reg [24:0] p6_add_35677;
  reg [24:0] p6_add_35678;
  reg [18:0] p6_add_35715;
  reg [18:0] p6_add_35718;
  reg [18:0] p6_add_35721;
  reg [18:0] p6_add_35724;
  reg [24:0] p6_add_35727;
  reg [24:0] p6_add_35728;
  reg [24:0] p6_add_35729;
  reg [24:0] p6_add_35730;
  reg [31:0] p6_umul_35592;
  reg [31:0] p6_umul_35598;
  reg [31:0] p6_umul_35604;
  reg [31:0] p6_umul_35610;
  reg [31:0] p6_umul_34389;
  reg [31:0] p6_umul_35622;
  reg [31:0] p6_umul_35623;
  reg [31:0] p6_umul_35624;
  reg [31:0] p6_umul_35626;
  reg [31:0] p6_umul_35627;
  reg [31:0] p6_umul_35628;
  reg [31:0] p6_umul_35630;
  reg [31:0] p6_umul_35631;
  reg [31:0] p6_umul_35632;
  reg [31:0] p6_umul_35634;
  reg [31:0] p6_umul_35635;
  reg [31:0] p6_umul_35636;
  reg [31:0] p6_umul_34412;
  reg [31:0] p6_umul_34413;
  reg [31:0] p6_umul_34416;
  always_ff @ (posedge clk) begin
    p6_bit_slice_35572 <= p6_bit_slice_35572_comb;
    p6_bit_slice_35576 <= p6_bit_slice_35576_comb;
    p6_bit_slice_35580 <= p6_bit_slice_35580_comb;
    p6_bit_slice_35584 <= p6_bit_slice_35584_comb;
    p6_bit_slice_35595 <= p6_bit_slice_35595_comb;
    p6_bit_slice_35601 <= p6_bit_slice_35601_comb;
    p6_bit_slice_35607 <= p6_bit_slice_35607_comb;
    p6_bit_slice_35613 <= p6_bit_slice_35613_comb;
    p6_bit_slice_35621 <= p6_bit_slice_35621_comb;
    p6_bit_slice_35625 <= p6_bit_slice_35625_comb;
    p6_bit_slice_35629 <= p6_bit_slice_35629_comb;
    p6_bit_slice_35633 <= p6_bit_slice_35633_comb;
    p6_bit_slice_35130 <= p5_bit_slice_35130;
    p6_bit_slice_35131 <= p5_bit_slice_35131;
    p6_bit_slice_35132 <= p5_bit_slice_35132;
    p6_bit_slice_35133 <= p5_bit_slice_35133;
    p6_bit_slice_35134 <= p5_bit_slice_35134;
    p6_bit_slice_35135 <= p5_bit_slice_35135;
    p6_bit_slice_35136 <= p5_bit_slice_35136;
    p6_bit_slice_35137 <= p5_bit_slice_35137;
    p6_bit_slice_33029 <= p5_bit_slice_33029;
    p6_bit_slice_33030 <= p5_bit_slice_33030;
    p6_bit_slice_33033 <= p5_bit_slice_33033;
    p6_bit_slice_33034 <= p5_bit_slice_33034;
    p6_sub_35679 <= p6_sub_35679_comb;
    p6_sub_35681 <= p6_sub_35681_comb;
    p6_sub_35683 <= p6_sub_35683_comb;
    p6_sub_35685 <= p6_sub_35685_comb;
    p6_bit_slice_35716 <= p6_bit_slice_35716_comb;
    p6_bit_slice_35717 <= p6_bit_slice_35717_comb;
    p6_bit_slice_35719 <= p6_bit_slice_35719_comb;
    p6_bit_slice_35720 <= p6_bit_slice_35720_comb;
    p6_bit_slice_35722 <= p6_bit_slice_35722_comb;
    p6_bit_slice_35723 <= p6_bit_slice_35723_comb;
    p6_bit_slice_35725 <= p6_bit_slice_35725_comb;
    p6_bit_slice_35726 <= p6_bit_slice_35726_comb;
    p6_bit_slice_35767 <= p6_bit_slice_35767_comb;
    p6_bit_slice_35768 <= p6_bit_slice_35768_comb;
    p6_bit_slice_35769 <= p6_bit_slice_35769_comb;
    p6_bit_slice_35770 <= p6_bit_slice_35770_comb;
    p6_bit_slice_35831 <= p6_bit_slice_35831_comb;
    p6_bit_slice_35832 <= p6_bit_slice_35832_comb;
    p6_bit_slice_35833 <= p6_bit_slice_35833_comb;
    p6_bit_slice_35834 <= p6_bit_slice_35834_comb;
    p6_bit_slice_35835 <= p6_bit_slice_35835_comb;
    p6_bit_slice_35836 <= p6_bit_slice_35836_comb;
    p6_bit_slice_35837 <= p6_bit_slice_35837_comb;
    p6_bit_slice_35838 <= p6_bit_slice_35838_comb;
    p6_bit_slice_35839 <= p6_bit_slice_35839_comb;
    p6_bit_slice_35840 <= p6_bit_slice_35840_comb;
    p6_bit_slice_35841 <= p6_bit_slice_35841_comb;
    p6_bit_slice_35842 <= p6_bit_slice_35842_comb;
    p6_bit_slice_35843 <= p6_bit_slice_35843_comb;
    p6_bit_slice_35844 <= p6_bit_slice_35844_comb;
    p6_bit_slice_35845 <= p6_bit_slice_35845_comb;
    p6_bit_slice_35846 <= p6_bit_slice_35846_comb;
    p6_add_35615 <= p6_add_35615_comb;
    p6_add_35618 <= p6_add_35618_comb;
    p6_add_35637 <= p6_add_35637_comb;
    p6_add_35638 <= p6_add_35638_comb;
    p6_add_35675 <= p6_add_35675_comb;
    p6_add_35676 <= p6_add_35676_comb;
    p6_add_35677 <= p6_add_35677_comb;
    p6_add_35678 <= p6_add_35678_comb;
    p6_add_35715 <= p6_add_35715_comb;
    p6_add_35718 <= p6_add_35718_comb;
    p6_add_35721 <= p6_add_35721_comb;
    p6_add_35724 <= p6_add_35724_comb;
    p6_add_35727 <= p6_add_35727_comb;
    p6_add_35728 <= p6_add_35728_comb;
    p6_add_35729 <= p6_add_35729_comb;
    p6_add_35730 <= p6_add_35730_comb;
    p6_umul_35592 <= p6_umul_35592_comb;
    p6_umul_35598 <= p6_umul_35598_comb;
    p6_umul_35604 <= p6_umul_35604_comb;
    p6_umul_35610 <= p6_umul_35610_comb;
    p6_umul_34389 <= p5_umul_34389;
    p6_umul_35622 <= p6_umul_35622_comb;
    p6_umul_35623 <= p6_umul_35623_comb;
    p6_umul_35624 <= p6_umul_35624_comb;
    p6_umul_35626 <= p6_umul_35626_comb;
    p6_umul_35627 <= p6_umul_35627_comb;
    p6_umul_35628 <= p6_umul_35628_comb;
    p6_umul_35630 <= p6_umul_35630_comb;
    p6_umul_35631 <= p6_umul_35631_comb;
    p6_umul_35632 <= p6_umul_35632_comb;
    p6_umul_35634 <= p6_umul_35634_comb;
    p6_umul_35635 <= p6_umul_35635_comb;
    p6_umul_35636 <= p6_umul_35636_comb;
    p6_umul_34412 <= p5_umul_34412;
    p6_umul_34413 <= p5_umul_34413;
    p6_umul_34416 <= p5_umul_34416;
  end

  // ===== Pipe stage 7:
  wire [23:0] p7_bit_slice_36307_comb;
  wire [23:0] p7_bit_slice_36308_comb;
  wire [23:0] p7_bit_slice_36309_comb;
  wire [23:0] p7_bit_slice_36310_comb;
  wire [28:0] p7_bit_slice_36311_comb;
  wire [28:0] p7_bit_slice_36312_comb;
  wire [28:0] p7_bit_slice_36313_comb;
  wire [28:0] p7_bit_slice_36314_comb;
  wire [23:0] p7_bit_slice_36051_comb;
  wire [23:0] p7_bit_slice_36052_comb;
  wire [23:0] p7_bit_slice_36070_comb;
  wire [23:0] p7_bit_slice_36072_comb;
  wire [31:0] p7_sign_ext_36323_comb;
  wire [31:0] p7_sign_ext_36324_comb;
  wire [31:0] p7_sign_ext_36325_comb;
  wire [31:0] p7_sign_ext_36326_comb;
  wire [31:0] p7_sign_ext_36327_comb;
  wire [31:0] p7_sign_ext_36328_comb;
  wire [31:0] p7_sign_ext_36329_comb;
  wire [31:0] p7_sign_ext_36330_comb;
  wire [29:0] p7_add_36036_comb;
  wire [29:0] p7_add_36038_comb;
  wire [29:0] p7_add_36040_comb;
  wire [29:0] p7_add_36042_comb;
  wire [31:0] p7_sign_ext_36069_comb;
  wire [31:0] p7_sign_ext_36071_comb;
  wire [31:0] p7_sign_ext_36100_comb;
  wire [31:0] p7_sign_ext_36104_comb;
  wire [31:0] p7_concat_36331_comb;
  wire [31:0] p7_concat_36333_comb;
  wire [31:0] p7_concat_36335_comb;
  wire [31:0] p7_concat_36337_comb;
  wire [23:0] p7_bit_slice_36349_comb;
  wire [23:0] p7_bit_slice_36352_comb;
  wire [23:0] p7_bit_slice_36355_comb;
  wire [23:0] p7_bit_slice_36358_comb;
  wire [31:0] p7_or_36043_comb;
  wire [31:0] p7_or_36045_comb;
  wire [31:0] p7_or_36047_comb;
  wire [31:0] p7_or_36049_comb;
  wire [31:0] p7_sub_36359_comb;
  wire [31:0] p7_sub_36360_comb;
  wire [31:0] p7_sub_36361_comb;
  wire [31:0] p7_sub_36362_comb;
  wire [18:0] p7_add_36363_comb;
  wire [18:0] p7_add_36365_comb;
  wire [18:0] p7_add_36367_comb;
  wire [18:0] p7_add_36369_comb;
  wire [31:0] p7_add_36371_comb;
  wire [31:0] p7_add_36372_comb;
  wire [31:0] p7_add_36373_comb;
  wire [31:0] p7_add_36374_comb;
  wire [18:0] p7_add_36375_comb;
  wire [31:0] p7_sign_ext_36377_comb;
  wire [18:0] p7_add_36378_comb;
  wire [31:0] p7_sign_ext_36380_comb;
  wire [18:0] p7_add_36381_comb;
  wire [31:0] p7_sign_ext_36383_comb;
  wire [18:0] p7_add_36384_comb;
  wire [31:0] p7_sign_ext_36386_comb;
  wire [29:0] p7_add_36053_comb;
  wire [31:0] p7_sub_36054_comb;
  wire [31:0] p7_sub_36055_comb;
  wire [31:0] p7_sub_36056_comb;
  wire [29:0] p7_add_36057_comb;
  wire [31:0] p7_sub_36058_comb;
  wire [31:0] p7_sub_36059_comb;
  wire [31:0] p7_sub_36060_comb;
  wire [29:0] p7_add_36061_comb;
  wire [31:0] p7_sub_36062_comb;
  wire [31:0] p7_sub_36063_comb;
  wire [31:0] p7_sub_36064_comb;
  wire [29:0] p7_add_36065_comb;
  wire [31:0] p7_sub_36066_comb;
  wire [31:0] p7_sub_36067_comb;
  wire [31:0] p7_sub_36068_comb;
  wire [24:0] p7_add_36137_comb;
  wire [20:0] p7_add_36139_comb;
  wire [24:0] p7_add_36144_comb;
  wire [20:0] p7_add_36146_comb;
  wire [24:0] p7_add_36151_comb;
  wire [29:0] p7_add_36152_comb;
  wire [24:0] p7_add_36157_comb;
  wire [28:0] p7_add_36158_comb;
  wire [24:0] p7_add_36177_comb;
  wire [20:0] p7_add_36179_comb;
  wire [24:0] p7_add_36183_comb;
  wire [20:0] p7_add_36185_comb;
  wire [24:0] p7_add_36189_comb;
  wire [29:0] p7_add_36190_comb;
  wire [24:0] p7_add_36193_comb;
  wire [28:0] p7_add_36194_comb;
  wire [28:0] p7_bit_slice_36073_comb;
  wire [28:0] p7_bit_slice_36074_comb;
  wire [28:0] p7_bit_slice_36075_comb;
  wire [28:0] p7_bit_slice_36076_comb;
  wire [28:0] p7_bit_slice_36077_comb;
  wire [28:0] p7_bit_slice_36078_comb;
  wire [28:0] p7_bit_slice_36079_comb;
  wire [28:0] p7_bit_slice_36080_comb;
  wire [28:0] p7_bit_slice_36081_comb;
  wire [28:0] p7_bit_slice_36082_comb;
  wire [28:0] p7_bit_slice_36083_comb;
  wire [28:0] p7_bit_slice_36084_comb;
  wire [28:0] p7_bit_slice_36085_comb;
  wire [28:0] p7_bit_slice_36086_comb;
  wire [28:0] p7_bit_slice_36087_comb;
  wire [28:0] p7_bit_slice_36088_comb;
  wire [31:0] p7_sign_ext_36089_comb;
  wire [31:0] p7_sign_ext_36090_comb;
  wire [31:0] p7_sign_ext_36091_comb;
  wire [31:0] p7_sign_ext_36092_comb;
  wire [31:0] p7_sign_ext_36093_comb;
  wire [31:0] p7_sign_ext_36094_comb;
  wire [31:0] p7_sign_ext_36095_comb;
  wire [31:0] p7_sign_ext_36096_comb;
  wire [23:0] p7_add_36411_comb;
  wire [23:0] p7_add_36413_comb;
  wire [23:0] p7_add_36415_comb;
  wire [23:0] p7_add_36417_comb;
  wire [23:0] p7_add_36419_comb;
  wire [23:0] p7_add_36421_comb;
  wire [23:0] p7_add_36422_comb;
  wire [23:0] p7_add_36424_comb;
  wire [23:0] p7_add_36425_comb;
  wire [23:0] p7_add_36427_comb;
  wire [23:0] p7_add_36428_comb;
  wire [23:0] p7_add_36430_comb;
  wire [23:0] p7_add_36435_comb;
  wire [23:0] p7_add_36437_comb;
  wire [23:0] p7_add_36439_comb;
  wire [23:0] p7_add_36441_comb;
  wire [23:0] p7_add_36443_comb;
  wire [23:0] p7_add_36444_comb;
  wire [23:0] p7_add_36446_comb;
  wire [23:0] p7_add_36447_comb;
  wire [23:0] p7_add_36449_comb;
  wire [23:0] p7_add_36450_comb;
  wire [23:0] p7_add_36452_comb;
  wire [23:0] p7_add_36453_comb;
  wire [31:0] p7_sign_ext_36113_comb;
  wire [31:0] p7_sign_ext_36114_comb;
  wire [31:0] p7_sign_ext_36115_comb;
  wire [31:0] p7_sign_ext_36116_comb;
  wire [31:0] p7_sign_ext_36117_comb;
  wire [31:0] p7_sign_ext_36118_comb;
  wire [31:0] p7_sign_ext_36119_comb;
  wire [31:0] p7_sign_ext_36120_comb;
  wire [31:0] p7_sign_ext_36121_comb;
  wire [31:0] p7_sign_ext_36122_comb;
  wire [31:0] p7_sign_ext_36123_comb;
  wire [31:0] p7_sign_ext_36124_comb;
  wire [31:0] p7_sign_ext_36125_comb;
  wire [31:0] p7_sign_ext_36126_comb;
  wire [31:0] p7_sign_ext_36127_comb;
  wire [31:0] p7_sign_ext_36128_comb;
  wire [31:0] p7_add_36129_comb;
  wire [31:0] p7_add_36131_comb;
  wire [31:0] p7_add_36133_comb;
  wire [31:0] p7_add_36135_comb;
  wire [29:0] p7_add_36203_comb;
  wire [20:0] p7_add_36205_comb;
  wire [28:0] p7_add_36209_comb;
  wire [20:0] p7_add_36211_comb;
  wire [20:0] p7_add_36215_comb;
  wire [20:0] p7_add_36218_comb;
  wire [20:0] p7_add_36223_comb;
  wire [20:0] p7_add_36226_comb;
  wire [29:0] p7_add_36249_comb;
  wire [20:0] p7_add_36251_comb;
  wire [28:0] p7_add_36255_comb;
  wire [20:0] p7_add_36257_comb;
  wire [20:0] p7_add_36261_comb;
  wire [20:0] p7_add_36264_comb;
  wire [20:0] p7_add_36269_comb;
  wire [20:0] p7_add_36272_comb;
  wire [31:0] p7_add_36163_comb;
  wire [31:0] p7_add_36164_comb;
  wire [31:0] p7_add_36165_comb;
  wire [31:0] p7_add_36166_comb;
  wire [31:0] p7_add_36167_comb;
  wire [31:0] p7_add_36168_comb;
  wire [31:0] p7_add_36169_comb;
  wire [31:0] p7_add_36170_comb;
  wire [31:0] p7_umul_36171_comb;
  wire [31:0] p7_umul_36172_comb;
  wire [31:0] p7_umul_36173_comb;
  wire [31:0] p7_umul_36174_comb;
  wire [31:0] p7_add_36232_comb;
  wire [31:0] p7_add_36233_comb;
  wire [31:0] p7_add_36235_comb;
  wire [31:0] p7_add_36236_comb;
  wire [31:0] p7_add_36238_comb;
  wire [31:0] p7_add_36239_comb;
  wire [31:0] p7_add_36241_comb;
  wire [31:0] p7_add_36242_comb;
  wire [31:0] p7_umul_36283_comb;
  wire [31:0] p7_umul_36284_comb;
  wire [31:0] p7_umul_36285_comb;
  wire [31:0] p7_umul_36286_comb;
  wire [31:0] p7_add_36483_comb;
  wire [31:0] p7_add_36484_comb;
  wire [31:0] p7_add_36485_comb;
  wire [31:0] p7_add_36486_comb;
  wire [31:0] p7_sub_36487_comb;
  wire [31:0] p7_sub_36488_comb;
  wire [31:0] p7_sub_36489_comb;
  wire [31:0] p7_sub_36490_comb;
  wire [31:0] p7_sub_36491_comb;
  wire [31:0] p7_sub_36492_comb;
  wire [31:0] p7_sub_36493_comb;
  wire [31:0] p7_sub_36494_comb;
  wire [31:0] p7_sub_36495_comb;
  wire [31:0] p7_sub_36496_comb;
  wire [31:0] p7_sub_36497_comb;
  wire [31:0] p7_sub_36498_comb;
  wire [31:0] p7_sub_36195_comb;
  wire [31:0] p7_sub_36196_comb;
  wire [31:0] p7_sub_36197_comb;
  wire [31:0] p7_sub_36198_comb;
  wire [29:0] p7_bit_slice_36199_comb;
  wire [29:0] p7_bit_slice_36200_comb;
  wire [29:0] p7_bit_slice_36201_comb;
  wire [29:0] p7_bit_slice_36202_comb;
  wire [31:0] p7_sub_36276_comb;
  wire [31:0] p7_sub_36278_comb;
  wire [31:0] p7_sub_36280_comb;
  wire [31:0] p7_sub_36282_comb;
  wire [31:0] p7_sub_36287_comb;
  wire [31:0] p7_sub_36290_comb;
  wire [31:0] p7_sub_36293_comb;
  wire [31:0] p7_sub_36296_comb;
  wire [26:0] p7_bit_slice_36299_comb;
  wire [26:0] p7_bit_slice_36300_comb;
  wire [26:0] p7_bit_slice_36301_comb;
  wire [26:0] p7_bit_slice_36302_comb;
  wire [31:0] p7_sub_36303_comb;
  wire [31:0] p7_sub_36304_comb;
  wire [31:0] p7_sub_36305_comb;
  wire [31:0] p7_sub_36306_comb;
  wire [31:0] p7_add_36431_comb;
  wire [31:0] p7_add_36432_comb;
  wire [31:0] p7_add_36433_comb;
  wire [31:0] p7_add_36434_comb;
  wire [31:0] p7_add_36455_comb;
  wire [31:0] p7_add_36456_comb;
  wire [31:0] p7_add_36457_comb;
  wire [31:0] p7_add_36458_comb;
  wire [17:0] p7_bit_slice_36499_comb;
  wire [17:0] p7_bit_slice_36500_comb;
  wire [17:0] p7_bit_slice_36501_comb;
  wire [17:0] p7_bit_slice_36502_comb;
  wire [17:0] p7_bit_slice_36503_comb;
  wire [17:0] p7_bit_slice_36504_comb;
  wire [17:0] p7_bit_slice_36505_comb;
  wire [17:0] p7_bit_slice_36506_comb;
  wire [17:0] p7_bit_slice_36507_comb;
  wire [17:0] p7_bit_slice_36508_comb;
  wire [17:0] p7_bit_slice_36509_comb;
  wire [17:0] p7_bit_slice_36510_comb;
  wire [17:0] p7_bit_slice_36511_comb;
  wire [17:0] p7_bit_slice_36512_comb;
  wire [17:0] p7_bit_slice_36513_comb;
  wire [17:0] p7_bit_slice_36514_comb;
  wire [31:0] p7_umul_36275_comb;
  wire [31:0] p7_umul_36277_comb;
  wire [31:0] p7_umul_36279_comb;
  wire [31:0] p7_umul_36281_comb;
  assign p7_bit_slice_36307_comb = p6_add_35675[24:1];
  assign p7_bit_slice_36308_comb = p6_add_35676[24:1];
  assign p7_bit_slice_36309_comb = p6_add_35677[24:1];
  assign p7_bit_slice_36310_comb = p6_add_35678[24:1];
  assign p7_bit_slice_36311_comb = p6_sub_35679[31:3];
  assign p7_bit_slice_36312_comb = p6_sub_35681[31:3];
  assign p7_bit_slice_36313_comb = p6_sub_35683[31:3];
  assign p7_bit_slice_36314_comb = p6_sub_35685[31:3];
  assign p7_bit_slice_36051_comb = p6_add_35615[24:1];
  assign p7_bit_slice_36052_comb = p6_add_35618[24:1];
  assign p7_bit_slice_36070_comb = p6_add_35637[24:1];
  assign p7_bit_slice_36072_comb = p6_add_35638[24:1];
  assign p7_sign_ext_36323_comb = {{8{p7_bit_slice_36307_comb[23]}}, p7_bit_slice_36307_comb};
  assign p7_sign_ext_36324_comb = {{8{p7_bit_slice_36308_comb[23]}}, p7_bit_slice_36308_comb};
  assign p7_sign_ext_36325_comb = {{8{p7_bit_slice_36309_comb[23]}}, p7_bit_slice_36309_comb};
  assign p7_sign_ext_36326_comb = {{8{p7_bit_slice_36310_comb[23]}}, p7_bit_slice_36310_comb};
  assign p7_sign_ext_36327_comb = {{3{p7_bit_slice_36311_comb[28]}}, p7_bit_slice_36311_comb};
  assign p7_sign_ext_36328_comb = {{3{p7_bit_slice_36312_comb[28]}}, p7_bit_slice_36312_comb};
  assign p7_sign_ext_36329_comb = {{3{p7_bit_slice_36313_comb[28]}}, p7_bit_slice_36313_comb};
  assign p7_sign_ext_36330_comb = {{3{p7_bit_slice_36314_comb[28]}}, p7_bit_slice_36314_comb};
  assign p7_add_36036_comb = p6_bit_slice_35572 + 30'h0000_0001;
  assign p7_add_36038_comb = p6_bit_slice_35576 + 30'h0000_0001;
  assign p7_add_36040_comb = p6_bit_slice_35580 + 30'h0000_0001;
  assign p7_add_36042_comb = p6_bit_slice_35584 + 30'h0000_0001;
  assign p7_sign_ext_36069_comb = {{8{p7_bit_slice_36051_comb[23]}}, p7_bit_slice_36051_comb};
  assign p7_sign_ext_36071_comb = {{8{p7_bit_slice_36052_comb[23]}}, p7_bit_slice_36052_comb};
  assign p7_sign_ext_36100_comb = {{8{p7_bit_slice_36070_comb[23]}}, p7_bit_slice_36070_comb};
  assign p7_sign_ext_36104_comb = {{8{p7_bit_slice_36072_comb[23]}}, p7_bit_slice_36072_comb};
  assign p7_concat_36331_comb = {p6_add_35715, p6_bit_slice_35716, 8'h00};
  assign p7_concat_36333_comb = {p6_add_35718, p6_bit_slice_35719, 8'h00};
  assign p7_concat_36335_comb = {p6_add_35721, p6_bit_slice_35722, 8'h00};
  assign p7_concat_36337_comb = {p6_add_35724, p6_bit_slice_35725, 8'h00};
  assign p7_bit_slice_36349_comb = p6_add_35727[24:1];
  assign p7_bit_slice_36352_comb = p6_add_35728[24:1];
  assign p7_bit_slice_36355_comb = p6_add_35729[24:1];
  assign p7_bit_slice_36358_comb = p6_add_35730[24:1];
  assign p7_or_36043_comb = p6_umul_35592 | 32'h0000_0004;
  assign p7_or_36045_comb = p6_umul_35598 | 32'h0000_0004;
  assign p7_or_36047_comb = p6_umul_35604 | 32'h0000_0004;
  assign p7_or_36049_comb = p6_umul_35610 | 32'h0000_0004;
  assign p7_sub_36359_comb = p7_concat_36331_comb - {p6_bit_slice_35717, 8'h00};
  assign p7_sub_36360_comb = p7_concat_36333_comb - {p6_bit_slice_35720, 8'h00};
  assign p7_sub_36361_comb = p7_concat_36335_comb - {p6_bit_slice_35723, 8'h00};
  assign p7_sub_36362_comb = p7_concat_36337_comb - {p6_bit_slice_35726, 8'h00};
  assign p7_add_36363_comb = p7_sign_ext_36323_comb[31:13] + 19'h0_0001;
  assign p7_add_36365_comb = p7_sign_ext_36324_comb[31:13] + 19'h0_0001;
  assign p7_add_36367_comb = p7_sign_ext_36325_comb[31:13] + 19'h0_0001;
  assign p7_add_36369_comb = p7_sign_ext_36326_comb[31:13] + 19'h0_0001;
  assign p7_add_36371_comb = p7_sign_ext_36323_comb + p7_sign_ext_36327_comb;
  assign p7_add_36372_comb = p7_sign_ext_36324_comb + p7_sign_ext_36328_comb;
  assign p7_add_36373_comb = p7_sign_ext_36325_comb + p7_sign_ext_36329_comb;
  assign p7_add_36374_comb = p7_sign_ext_36326_comb + p7_sign_ext_36330_comb;
  assign p7_add_36375_comb = p7_sign_ext_36327_comb[31:13] + 19'h0_0001;
  assign p7_sign_ext_36377_comb = {{8{p7_bit_slice_36349_comb[23]}}, p7_bit_slice_36349_comb};
  assign p7_add_36378_comb = p7_sign_ext_36328_comb[31:13] + 19'h0_0001;
  assign p7_sign_ext_36380_comb = {{8{p7_bit_slice_36352_comb[23]}}, p7_bit_slice_36352_comb};
  assign p7_add_36381_comb = p7_sign_ext_36329_comb[31:13] + 19'h0_0001;
  assign p7_sign_ext_36383_comb = {{8{p7_bit_slice_36355_comb[23]}}, p7_bit_slice_36355_comb};
  assign p7_add_36384_comb = p7_sign_ext_36330_comb[31:13] + 19'h0_0001;
  assign p7_sign_ext_36386_comb = {{8{p7_bit_slice_36358_comb[23]}}, p7_bit_slice_36358_comb};
  assign p7_add_36053_comb = p6_bit_slice_35621 + p7_add_36036_comb;
  assign p7_sub_36054_comb = p7_or_36043_comb - p6_umul_35622;
  assign p7_sub_36055_comb = p7_or_36043_comb - p6_umul_35623;
  assign p7_sub_36056_comb = {p7_add_36036_comb, p6_bit_slice_35595} - p6_umul_35624;
  assign p7_add_36057_comb = p6_bit_slice_35625 + p7_add_36038_comb;
  assign p7_sub_36058_comb = p7_or_36045_comb - p6_umul_35626;
  assign p7_sub_36059_comb = p7_or_36045_comb - p6_umul_35627;
  assign p7_sub_36060_comb = {p7_add_36038_comb, p6_bit_slice_35601} - p6_umul_35628;
  assign p7_add_36061_comb = p6_bit_slice_35629 + p7_add_36040_comb;
  assign p7_sub_36062_comb = p7_or_36047_comb - p6_umul_35630;
  assign p7_sub_36063_comb = p7_or_36047_comb - p6_umul_35631;
  assign p7_sub_36064_comb = {p7_add_36040_comb, p6_bit_slice_35607} - p6_umul_35632;
  assign p7_add_36065_comb = p6_bit_slice_35633 + p7_add_36042_comb;
  assign p7_sub_36066_comb = p7_or_36049_comb - p6_umul_35634;
  assign p7_sub_36067_comb = p7_or_36049_comb - p6_umul_35635;
  assign p7_sub_36068_comb = {p7_add_36042_comb, p6_bit_slice_35613} - p6_umul_35636;
  assign p7_add_36137_comb = p7_sign_ext_36069_comb[31:7] + 25'h000_0001;
  assign p7_add_36139_comb = p6_umul_34389[31:11] + p6_bit_slice_33030;
  assign p7_add_36144_comb = p7_sign_ext_36071_comb[31:7] + 25'h000_0001;
  assign p7_add_36146_comb = p6_umul_34413[31:11] + p6_bit_slice_33030;
  assign p7_add_36151_comb = p6_umul_34413[31:7] + 25'h000_0001;
  assign p7_add_36152_comb = p7_sign_ext_36071_comb[31:2] + p6_umul_34389[31:2];
  assign p7_add_36157_comb = p6_umul_34389[31:7] + 25'h000_0001;
  assign p7_add_36158_comb = p7_sign_ext_36069_comb[31:3] + p6_umul_34413[31:3];
  assign p7_add_36177_comb = p7_sign_ext_36100_comb[31:7] + 25'h000_0001;
  assign p7_add_36179_comb = p6_umul_34412[31:11] + p6_bit_slice_33034;
  assign p7_add_36183_comb = p7_sign_ext_36104_comb[31:7] + 25'h000_0001;
  assign p7_add_36185_comb = p6_umul_34416[31:11] + p6_bit_slice_33034;
  assign p7_add_36189_comb = p6_umul_34416[31:7] + 25'h000_0001;
  assign p7_add_36190_comb = p7_sign_ext_36104_comb[31:2] + p6_umul_34412[31:2];
  assign p7_add_36193_comb = p6_umul_34412[31:7] + 25'h000_0001;
  assign p7_add_36194_comb = p7_sign_ext_36100_comb[31:3] + p6_umul_34416[31:3];
  assign p7_bit_slice_36073_comb = p7_add_36053_comb[29:1];
  assign p7_bit_slice_36074_comb = p7_sub_36054_comb[31:3];
  assign p7_bit_slice_36075_comb = p7_sub_36055_comb[31:3];
  assign p7_bit_slice_36076_comb = p7_sub_36056_comb[31:3];
  assign p7_bit_slice_36077_comb = p7_add_36057_comb[29:1];
  assign p7_bit_slice_36078_comb = p7_sub_36058_comb[31:3];
  assign p7_bit_slice_36079_comb = p7_sub_36059_comb[31:3];
  assign p7_bit_slice_36080_comb = p7_sub_36060_comb[31:3];
  assign p7_bit_slice_36081_comb = p7_add_36061_comb[29:1];
  assign p7_bit_slice_36082_comb = p7_sub_36062_comb[31:3];
  assign p7_bit_slice_36083_comb = p7_sub_36063_comb[31:3];
  assign p7_bit_slice_36084_comb = p7_sub_36064_comb[31:3];
  assign p7_bit_slice_36085_comb = p7_add_36065_comb[29:1];
  assign p7_bit_slice_36086_comb = p7_sub_36066_comb[31:3];
  assign p7_bit_slice_36087_comb = p7_sub_36067_comb[31:3];
  assign p7_bit_slice_36088_comb = p7_sub_36068_comb[31:3];
  assign p7_sign_ext_36089_comb = {{8{p6_bit_slice_35130[23]}}, p6_bit_slice_35130};
  assign p7_sign_ext_36090_comb = {{8{p6_bit_slice_35131[23]}}, p6_bit_slice_35131};
  assign p7_sign_ext_36091_comb = {{8{p6_bit_slice_35132[23]}}, p6_bit_slice_35132};
  assign p7_sign_ext_36092_comb = {{8{p6_bit_slice_35133[23]}}, p6_bit_slice_35133};
  assign p7_sign_ext_36093_comb = {{8{p6_bit_slice_35134[23]}}, p6_bit_slice_35134};
  assign p7_sign_ext_36094_comb = {{8{p6_bit_slice_35135[23]}}, p6_bit_slice_35135};
  assign p7_sign_ext_36095_comb = {{8{p6_bit_slice_35136[23]}}, p6_bit_slice_35136};
  assign p7_sign_ext_36096_comb = {{8{p6_bit_slice_35137[23]}}, p6_bit_slice_35137};
  assign p7_add_36411_comb = p7_sign_ext_36327_comb[31:8] + p7_sub_36359_comb[31:8];
  assign p7_add_36413_comb = p7_sign_ext_36328_comb[31:8] + p7_sub_36360_comb[31:8];
  assign p7_add_36415_comb = p7_sign_ext_36329_comb[31:8] + p7_sub_36361_comb[31:8];
  assign p7_add_36417_comb = p7_sign_ext_36330_comb[31:8] + p7_sub_36362_comb[31:8];
  assign p7_add_36419_comb = {p7_add_36363_comb, p6_add_35675[13:9]} + p6_bit_slice_35767;
  assign p7_add_36421_comb = p7_sign_ext_36327_comb[31:8] + p6_bit_slice_35717;
  assign p7_add_36422_comb = {p7_add_36365_comb, p6_add_35676[13:9]} + p6_bit_slice_35768;
  assign p7_add_36424_comb = p7_sign_ext_36328_comb[31:8] + p6_bit_slice_35720;
  assign p7_add_36425_comb = {p7_add_36367_comb, p6_add_35677[13:9]} + p6_bit_slice_35769;
  assign p7_add_36427_comb = p7_sign_ext_36329_comb[31:8] + p6_bit_slice_35723;
  assign p7_add_36428_comb = {p7_add_36369_comb, p6_add_35678[13:9]} + p6_bit_slice_35770;
  assign p7_add_36430_comb = p7_sign_ext_36330_comb[31:8] + p6_bit_slice_35726;
  assign p7_add_36435_comb = p7_add_36371_comb[31:8] + p6_bit_slice_35717;
  assign p7_add_36437_comb = p7_add_36372_comb[31:8] + p6_bit_slice_35720;
  assign p7_add_36439_comb = p7_add_36373_comb[31:8] + p6_bit_slice_35723;
  assign p7_add_36441_comb = p7_add_36374_comb[31:8] + p6_bit_slice_35726;
  assign p7_add_36443_comb = {p7_add_36375_comb, p6_sub_35679[15:11]} + p6_bit_slice_35767;
  assign p7_add_36444_comb = p7_sign_ext_36377_comb[31:8] + p6_bit_slice_35717;
  assign p7_add_36446_comb = {p7_add_36378_comb, p6_sub_35681[15:11]} + p6_bit_slice_35768;
  assign p7_add_36447_comb = p7_sign_ext_36380_comb[31:8] + p6_bit_slice_35720;
  assign p7_add_36449_comb = {p7_add_36381_comb, p6_sub_35683[15:11]} + p6_bit_slice_35769;
  assign p7_add_36450_comb = p7_sign_ext_36383_comb[31:8] + p6_bit_slice_35723;
  assign p7_add_36452_comb = {p7_add_36384_comb, p6_sub_35685[15:11]} + p6_bit_slice_35770;
  assign p7_add_36453_comb = p7_sign_ext_36386_comb[31:8] + p6_bit_slice_35726;
  assign p7_sign_ext_36113_comb = {{3{p7_bit_slice_36073_comb[28]}}, p7_bit_slice_36073_comb};
  assign p7_sign_ext_36114_comb = {{3{p7_bit_slice_36074_comb[28]}}, p7_bit_slice_36074_comb};
  assign p7_sign_ext_36115_comb = {{3{p7_bit_slice_36075_comb[28]}}, p7_bit_slice_36075_comb};
  assign p7_sign_ext_36116_comb = {{3{p7_bit_slice_36076_comb[28]}}, p7_bit_slice_36076_comb};
  assign p7_sign_ext_36117_comb = {{3{p7_bit_slice_36077_comb[28]}}, p7_bit_slice_36077_comb};
  assign p7_sign_ext_36118_comb = {{3{p7_bit_slice_36078_comb[28]}}, p7_bit_slice_36078_comb};
  assign p7_sign_ext_36119_comb = {{3{p7_bit_slice_36079_comb[28]}}, p7_bit_slice_36079_comb};
  assign p7_sign_ext_36120_comb = {{3{p7_bit_slice_36080_comb[28]}}, p7_bit_slice_36080_comb};
  assign p7_sign_ext_36121_comb = {{3{p7_bit_slice_36081_comb[28]}}, p7_bit_slice_36081_comb};
  assign p7_sign_ext_36122_comb = {{3{p7_bit_slice_36082_comb[28]}}, p7_bit_slice_36082_comb};
  assign p7_sign_ext_36123_comb = {{3{p7_bit_slice_36083_comb[28]}}, p7_bit_slice_36083_comb};
  assign p7_sign_ext_36124_comb = {{3{p7_bit_slice_36084_comb[28]}}, p7_bit_slice_36084_comb};
  assign p7_sign_ext_36125_comb = {{3{p7_bit_slice_36085_comb[28]}}, p7_bit_slice_36085_comb};
  assign p7_sign_ext_36126_comb = {{3{p7_bit_slice_36086_comb[28]}}, p7_bit_slice_36086_comb};
  assign p7_sign_ext_36127_comb = {{3{p7_bit_slice_36087_comb[28]}}, p7_bit_slice_36087_comb};
  assign p7_sign_ext_36128_comb = {{3{p7_bit_slice_36088_comb[28]}}, p7_bit_slice_36088_comb};
  assign p7_add_36129_comb = p7_sign_ext_36089_comb + p7_sign_ext_36090_comb;
  assign p7_add_36131_comb = p7_sign_ext_36091_comb + p7_sign_ext_36092_comb;
  assign p7_add_36133_comb = p7_sign_ext_36093_comb + p7_sign_ext_36094_comb;
  assign p7_add_36135_comb = p7_sign_ext_36095_comb + p7_sign_ext_36096_comb;
  assign p7_add_36203_comb = {p7_add_36137_comb, p6_add_35615[7:3]} + {p7_add_36139_comb, p6_umul_34389[10:2]};
  assign p7_add_36205_comb = p6_umul_34413[31:11] + p6_bit_slice_33029;
  assign p7_add_36209_comb = {p7_add_36144_comb, p6_add_35618[7:4]} + {p7_add_36146_comb, p6_umul_34413[10:3]};
  assign p7_add_36211_comb = p6_umul_34389[31:11] + p6_bit_slice_33029;
  assign p7_add_36215_comb = p7_add_36151_comb[24:4] + p6_bit_slice_33030;
  assign p7_add_36218_comb = p7_add_36152_comb[29:9] + p6_bit_slice_33029;
  assign p7_add_36223_comb = p7_add_36157_comb[24:4] + p6_bit_slice_33030;
  assign p7_add_36226_comb = p7_add_36158_comb[28:8] + p6_bit_slice_33029;
  assign p7_add_36249_comb = {p7_add_36177_comb, p6_add_35637[7:3]} + {p7_add_36179_comb, p6_umul_34412[10:2]};
  assign p7_add_36251_comb = p6_umul_34416[31:11] + p6_bit_slice_33033;
  assign p7_add_36255_comb = {p7_add_36183_comb, p6_add_35638[7:4]} + {p7_add_36185_comb, p6_umul_34416[10:3]};
  assign p7_add_36257_comb = p6_umul_34412[31:11] + p6_bit_slice_33033;
  assign p7_add_36261_comb = p7_add_36189_comb[24:4] + p6_bit_slice_33034;
  assign p7_add_36264_comb = p7_add_36190_comb[29:9] + p6_bit_slice_33033;
  assign p7_add_36269_comb = p7_add_36193_comb[24:4] + p6_bit_slice_33034;
  assign p7_add_36272_comb = p7_add_36194_comb[28:8] + p6_bit_slice_33033;
  assign p7_add_36163_comb = p7_sign_ext_36113_comb + p7_sign_ext_36114_comb;
  assign p7_add_36164_comb = p7_sign_ext_36115_comb + p7_sign_ext_36116_comb;
  assign p7_add_36165_comb = p7_sign_ext_36117_comb + p7_sign_ext_36118_comb;
  assign p7_add_36166_comb = p7_sign_ext_36119_comb + p7_sign_ext_36120_comb;
  assign p7_add_36167_comb = p7_sign_ext_36121_comb + p7_sign_ext_36122_comb;
  assign p7_add_36168_comb = p7_sign_ext_36123_comb + p7_sign_ext_36124_comb;
  assign p7_add_36169_comb = p7_sign_ext_36125_comb + p7_sign_ext_36126_comb;
  assign p7_add_36170_comb = p7_sign_ext_36127_comb + p7_sign_ext_36128_comb;
  assign p7_umul_36171_comb = umul32b_32b_x_11b(p7_add_36129_comb, 11'h454);
  assign p7_umul_36172_comb = umul32b_32b_x_11b(p7_add_36131_comb, 11'h454);
  assign p7_umul_36173_comb = umul32b_32b_x_11b(p7_add_36133_comb, 11'h454);
  assign p7_umul_36174_comb = umul32b_32b_x_11b(p7_add_36135_comb, 11'h454);
  assign p7_add_36232_comb = p7_sign_ext_36113_comb + p7_sign_ext_36116_comb;
  assign p7_add_36233_comb = p7_sign_ext_36115_comb + p7_sign_ext_36114_comb;
  assign p7_add_36235_comb = p7_sign_ext_36117_comb + p7_sign_ext_36120_comb;
  assign p7_add_36236_comb = p7_sign_ext_36119_comb + p7_sign_ext_36118_comb;
  assign p7_add_36238_comb = p7_sign_ext_36121_comb + p7_sign_ext_36124_comb;
  assign p7_add_36239_comb = p7_sign_ext_36123_comb + p7_sign_ext_36122_comb;
  assign p7_add_36241_comb = p7_sign_ext_36125_comb + p7_sign_ext_36128_comb;
  assign p7_add_36242_comb = p7_sign_ext_36127_comb + p7_sign_ext_36126_comb;
  assign p7_umul_36283_comb = umul32b_32b_x_11b(p7_sign_ext_36089_comb, 11'h620);
  assign p7_umul_36284_comb = umul32b_32b_x_11b(p7_sign_ext_36091_comb, 11'h620);
  assign p7_umul_36285_comb = umul32b_32b_x_11b(p7_sign_ext_36093_comb, 11'h620);
  assign p7_umul_36286_comb = umul32b_32b_x_11b(p7_sign_ext_36095_comb, 11'h620);
  assign p7_add_36483_comb = p7_sign_ext_36377_comb + {p7_add_36411_comb, p6_sub_35679[10:3]};
  assign p7_add_36484_comb = p7_sign_ext_36380_comb + {p7_add_36413_comb, p6_sub_35681[10:3]};
  assign p7_add_36485_comb = p7_sign_ext_36383_comb + {p7_add_36415_comb, p6_sub_35683[10:3]};
  assign p7_add_36486_comb = p7_sign_ext_36386_comb + {p7_add_36417_comb, p6_sub_35685[10:3]};
  assign p7_sub_36487_comb = {p7_add_36419_comb, p6_add_35675[8:1]} - {p7_add_36421_comb, p6_sub_35679[10:3]};
  assign p7_sub_36488_comb = {p7_add_36422_comb, p6_add_35676[8:1]} - {p7_add_36424_comb, p6_sub_35681[10:3]};
  assign p7_sub_36489_comb = {p7_add_36425_comb, p6_add_35677[8:1]} - {p7_add_36427_comb, p6_sub_35683[10:3]};
  assign p7_sub_36490_comb = {p7_add_36428_comb, p6_add_35678[8:1]} - {p7_add_36430_comb, p6_sub_35685[10:3]};
  assign p7_sub_36491_comb = p7_concat_36331_comb - {p7_add_36435_comb, p7_add_36371_comb[7:0]};
  assign p7_sub_36492_comb = p7_concat_36333_comb - {p7_add_36437_comb, p7_add_36372_comb[7:0]};
  assign p7_sub_36493_comb = p7_concat_36335_comb - {p7_add_36439_comb, p7_add_36373_comb[7:0]};
  assign p7_sub_36494_comb = p7_concat_36337_comb - {p7_add_36441_comb, p7_add_36374_comb[7:0]};
  assign p7_sub_36495_comb = {p7_add_36443_comb, p6_sub_35679[10:3]} - {p7_add_36444_comb, p6_add_35727[8:1]};
  assign p7_sub_36496_comb = {p7_add_36446_comb, p6_sub_35681[10:3]} - {p7_add_36447_comb, p6_add_35728[8:1]};
  assign p7_sub_36497_comb = {p7_add_36449_comb, p6_sub_35683[10:3]} - {p7_add_36450_comb, p6_add_35729[8:1]};
  assign p7_sub_36498_comb = {p7_add_36452_comb, p6_sub_35685[10:3]} - {p7_add_36453_comb, p6_add_35730[8:1]};
  assign p7_sub_36195_comb = p7_add_36163_comb - p7_add_36164_comb;
  assign p7_sub_36196_comb = p7_add_36165_comb - p7_add_36166_comb;
  assign p7_sub_36197_comb = p7_add_36167_comb - p7_add_36168_comb;
  assign p7_sub_36198_comb = p7_add_36169_comb - p7_add_36170_comb;
  assign p7_bit_slice_36199_comb = p7_umul_36171_comb[31:2];
  assign p7_bit_slice_36200_comb = p7_umul_36172_comb[31:2];
  assign p7_bit_slice_36201_comb = p7_umul_36173_comb[31:2];
  assign p7_bit_slice_36202_comb = p7_umul_36174_comb[31:2];
  assign p7_sub_36276_comb = p7_add_36232_comb - p7_add_36233_comb;
  assign p7_sub_36278_comb = p7_add_36235_comb - p7_add_36236_comb;
  assign p7_sub_36280_comb = p7_add_36238_comb - p7_add_36239_comb;
  assign p7_sub_36282_comb = p7_add_36241_comb - p7_add_36242_comb;
  assign p7_sub_36287_comb = {p7_add_36203_comb, p6_add_35615[2:1]} - {p7_add_36205_comb, p6_umul_34413[10:0]};
  assign p7_sub_36290_comb = {p7_add_36209_comb, p6_add_35618[3:1]} - {p7_add_36211_comb, p6_umul_34389[10:0]};
  assign p7_sub_36293_comb = {p7_add_36215_comb, p7_add_36151_comb[3:0], p6_umul_34413[6:0]} - {p7_add_36218_comb, p7_add_36152_comb[8:0], p6_add_35618[2:1]};
  assign p7_sub_36296_comb = {p7_add_36223_comb, p7_add_36157_comb[3:0], p6_umul_34389[6:0]} - {p7_add_36226_comb, p7_add_36158_comb[7:0], p6_add_35615[3:1]};
  assign p7_bit_slice_36299_comb = p7_umul_36283_comb[31:5];
  assign p7_bit_slice_36300_comb = p7_umul_36284_comb[31:5];
  assign p7_bit_slice_36301_comb = p7_umul_36285_comb[31:5];
  assign p7_bit_slice_36302_comb = p7_umul_36286_comb[31:5];
  assign p7_sub_36303_comb = {p7_add_36249_comb, p6_add_35637[2:1]} - {p7_add_36251_comb, p6_umul_34416[10:0]};
  assign p7_sub_36304_comb = {p7_add_36255_comb, p6_add_35638[3:1]} - {p7_add_36257_comb, p6_umul_34412[10:0]};
  assign p7_sub_36305_comb = {p7_add_36261_comb, p7_add_36189_comb[3:0], p6_umul_34416[6:0]} - {p7_add_36264_comb, p7_add_36190_comb[8:0], p6_add_35638[2:1]};
  assign p7_sub_36306_comb = {p7_add_36269_comb, p7_add_36193_comb[3:0], p6_umul_34412[6:0]} - {p7_add_36272_comb, p7_add_36194_comb[7:0], p6_add_35637[3:1]};
  assign p7_add_36431_comb = p7_sign_ext_36114_comb + p7_sign_ext_36116_comb;
  assign p7_add_36432_comb = p7_sign_ext_36118_comb + p7_sign_ext_36120_comb;
  assign p7_add_36433_comb = p7_sign_ext_36122_comb + p7_sign_ext_36124_comb;
  assign p7_add_36434_comb = p7_sign_ext_36126_comb + p7_sign_ext_36128_comb;
  assign p7_add_36455_comb = p7_sign_ext_36115_comb + p7_sign_ext_36113_comb;
  assign p7_add_36456_comb = p7_sign_ext_36119_comb + p7_sign_ext_36117_comb;
  assign p7_add_36457_comb = p7_sign_ext_36123_comb + p7_sign_ext_36121_comb;
  assign p7_add_36458_comb = p7_sign_ext_36127_comb + p7_sign_ext_36125_comb;
  assign p7_bit_slice_36499_comb = p7_add_36483_comb[31:14];
  assign p7_bit_slice_36500_comb = p7_add_36484_comb[31:14];
  assign p7_bit_slice_36501_comb = p7_add_36485_comb[31:14];
  assign p7_bit_slice_36502_comb = p7_add_36486_comb[31:14];
  assign p7_bit_slice_36503_comb = p7_sub_36487_comb[31:14];
  assign p7_bit_slice_36504_comb = p7_sub_36488_comb[31:14];
  assign p7_bit_slice_36505_comb = p7_sub_36489_comb[31:14];
  assign p7_bit_slice_36506_comb = p7_sub_36490_comb[31:14];
  assign p7_bit_slice_36507_comb = p7_sub_36491_comb[31:14];
  assign p7_bit_slice_36508_comb = p7_sub_36492_comb[31:14];
  assign p7_bit_slice_36509_comb = p7_sub_36493_comb[31:14];
  assign p7_bit_slice_36510_comb = p7_sub_36494_comb[31:14];
  assign p7_bit_slice_36511_comb = p7_sub_36495_comb[31:14];
  assign p7_bit_slice_36512_comb = p7_sub_36496_comb[31:14];
  assign p7_bit_slice_36513_comb = p7_sub_36497_comb[31:14];
  assign p7_bit_slice_36514_comb = p7_sub_36498_comb[31:14];
  assign p7_umul_36275_comb = umul32b_32b_x_12b(p7_sign_ext_36090_comb, 12'hec8);
  assign p7_umul_36277_comb = umul32b_32b_x_12b(p7_sign_ext_36092_comb, 12'hec8);
  assign p7_umul_36279_comb = umul32b_32b_x_12b(p7_sign_ext_36094_comb, 12'hec8);
  assign p7_umul_36281_comb = umul32b_32b_x_12b(p7_sign_ext_36096_comb, 12'hec8);

  // Registers for pipe stage 7:
  reg [31:0] p7_sub_36195;
  reg [31:0] p7_sub_36196;
  reg [31:0] p7_sub_36197;
  reg [31:0] p7_sub_36198;
  reg [29:0] p7_bit_slice_36199;
  reg [29:0] p7_bit_slice_36200;
  reg [29:0] p7_bit_slice_36201;
  reg [29:0] p7_bit_slice_36202;
  reg [31:0] p7_sub_36276;
  reg [31:0] p7_sub_36278;
  reg [31:0] p7_sub_36280;
  reg [31:0] p7_sub_36282;
  reg [31:0] p7_sub_36287;
  reg [31:0] p7_sub_36290;
  reg [31:0] p7_sub_36293;
  reg [31:0] p7_sub_36296;
  reg [26:0] p7_bit_slice_36299;
  reg [26:0] p7_bit_slice_36300;
  reg [26:0] p7_bit_slice_36301;
  reg [26:0] p7_bit_slice_36302;
  reg [31:0] p7_sub_36303;
  reg [31:0] p7_sub_36304;
  reg [31:0] p7_sub_36305;
  reg [31:0] p7_sub_36306;
  reg [31:0] p7_add_36431;
  reg [31:0] p7_add_36432;
  reg [31:0] p7_add_36433;
  reg [31:0] p7_add_36434;
  reg [31:0] p7_add_36455;
  reg [31:0] p7_add_36456;
  reg [31:0] p7_add_36457;
  reg [31:0] p7_add_36458;
  reg [17:0] p7_bit_slice_35831;
  reg [17:0] p7_bit_slice_35832;
  reg [17:0] p7_bit_slice_35833;
  reg [17:0] p7_bit_slice_35834;
  reg [17:0] p7_bit_slice_36499;
  reg [17:0] p7_bit_slice_36500;
  reg [17:0] p7_bit_slice_36501;
  reg [17:0] p7_bit_slice_36502;
  reg [17:0] p7_bit_slice_36503;
  reg [17:0] p7_bit_slice_36504;
  reg [17:0] p7_bit_slice_36505;
  reg [17:0] p7_bit_slice_36506;
  reg [17:0] p7_bit_slice_35835;
  reg [17:0] p7_bit_slice_35836;
  reg [17:0] p7_bit_slice_35837;
  reg [17:0] p7_bit_slice_35838;
  reg [17:0] p7_bit_slice_35839;
  reg [17:0] p7_bit_slice_35840;
  reg [17:0] p7_bit_slice_35841;
  reg [17:0] p7_bit_slice_35842;
  reg [17:0] p7_bit_slice_36507;
  reg [17:0] p7_bit_slice_36508;
  reg [17:0] p7_bit_slice_36509;
  reg [17:0] p7_bit_slice_36510;
  reg [17:0] p7_bit_slice_36511;
  reg [17:0] p7_bit_slice_36512;
  reg [17:0] p7_bit_slice_36513;
  reg [17:0] p7_bit_slice_36514;
  reg [17:0] p7_bit_slice_35843;
  reg [17:0] p7_bit_slice_35844;
  reg [17:0] p7_bit_slice_35845;
  reg [17:0] p7_bit_slice_35846;
  reg [31:0] p7_umul_36275;
  reg [31:0] p7_umul_36277;
  reg [31:0] p7_umul_36279;
  reg [31:0] p7_umul_36281;
  always_ff @ (posedge clk) begin
    p7_sub_36195 <= p7_sub_36195_comb;
    p7_sub_36196 <= p7_sub_36196_comb;
    p7_sub_36197 <= p7_sub_36197_comb;
    p7_sub_36198 <= p7_sub_36198_comb;
    p7_bit_slice_36199 <= p7_bit_slice_36199_comb;
    p7_bit_slice_36200 <= p7_bit_slice_36200_comb;
    p7_bit_slice_36201 <= p7_bit_slice_36201_comb;
    p7_bit_slice_36202 <= p7_bit_slice_36202_comb;
    p7_sub_36276 <= p7_sub_36276_comb;
    p7_sub_36278 <= p7_sub_36278_comb;
    p7_sub_36280 <= p7_sub_36280_comb;
    p7_sub_36282 <= p7_sub_36282_comb;
    p7_sub_36287 <= p7_sub_36287_comb;
    p7_sub_36290 <= p7_sub_36290_comb;
    p7_sub_36293 <= p7_sub_36293_comb;
    p7_sub_36296 <= p7_sub_36296_comb;
    p7_bit_slice_36299 <= p7_bit_slice_36299_comb;
    p7_bit_slice_36300 <= p7_bit_slice_36300_comb;
    p7_bit_slice_36301 <= p7_bit_slice_36301_comb;
    p7_bit_slice_36302 <= p7_bit_slice_36302_comb;
    p7_sub_36303 <= p7_sub_36303_comb;
    p7_sub_36304 <= p7_sub_36304_comb;
    p7_sub_36305 <= p7_sub_36305_comb;
    p7_sub_36306 <= p7_sub_36306_comb;
    p7_add_36431 <= p7_add_36431_comb;
    p7_add_36432 <= p7_add_36432_comb;
    p7_add_36433 <= p7_add_36433_comb;
    p7_add_36434 <= p7_add_36434_comb;
    p7_add_36455 <= p7_add_36455_comb;
    p7_add_36456 <= p7_add_36456_comb;
    p7_add_36457 <= p7_add_36457_comb;
    p7_add_36458 <= p7_add_36458_comb;
    p7_bit_slice_35831 <= p6_bit_slice_35831;
    p7_bit_slice_35832 <= p6_bit_slice_35832;
    p7_bit_slice_35833 <= p6_bit_slice_35833;
    p7_bit_slice_35834 <= p6_bit_slice_35834;
    p7_bit_slice_36499 <= p7_bit_slice_36499_comb;
    p7_bit_slice_36500 <= p7_bit_slice_36500_comb;
    p7_bit_slice_36501 <= p7_bit_slice_36501_comb;
    p7_bit_slice_36502 <= p7_bit_slice_36502_comb;
    p7_bit_slice_36503 <= p7_bit_slice_36503_comb;
    p7_bit_slice_36504 <= p7_bit_slice_36504_comb;
    p7_bit_slice_36505 <= p7_bit_slice_36505_comb;
    p7_bit_slice_36506 <= p7_bit_slice_36506_comb;
    p7_bit_slice_35835 <= p6_bit_slice_35835;
    p7_bit_slice_35836 <= p6_bit_slice_35836;
    p7_bit_slice_35837 <= p6_bit_slice_35837;
    p7_bit_slice_35838 <= p6_bit_slice_35838;
    p7_bit_slice_35839 <= p6_bit_slice_35839;
    p7_bit_slice_35840 <= p6_bit_slice_35840;
    p7_bit_slice_35841 <= p6_bit_slice_35841;
    p7_bit_slice_35842 <= p6_bit_slice_35842;
    p7_bit_slice_36507 <= p7_bit_slice_36507_comb;
    p7_bit_slice_36508 <= p7_bit_slice_36508_comb;
    p7_bit_slice_36509 <= p7_bit_slice_36509_comb;
    p7_bit_slice_36510 <= p7_bit_slice_36510_comb;
    p7_bit_slice_36511 <= p7_bit_slice_36511_comb;
    p7_bit_slice_36512 <= p7_bit_slice_36512_comb;
    p7_bit_slice_36513 <= p7_bit_slice_36513_comb;
    p7_bit_slice_36514 <= p7_bit_slice_36514_comb;
    p7_bit_slice_35843 <= p6_bit_slice_35843;
    p7_bit_slice_35844 <= p6_bit_slice_35844;
    p7_bit_slice_35845 <= p6_bit_slice_35845;
    p7_bit_slice_35846 <= p6_bit_slice_35846;
    p7_umul_36275 <= p7_umul_36275_comb;
    p7_umul_36277 <= p7_umul_36277_comb;
    p7_umul_36279 <= p7_umul_36279_comb;
    p7_umul_36281 <= p7_umul_36281_comb;
  end

  // ===== Pipe stage 8:
  wire [29:0] p8_add_36663_comb;
  wire [29:0] p8_add_36665_comb;
  wire [29:0] p8_add_36667_comb;
  wire [29:0] p8_add_36669_comb;
  wire [26:0] p8_add_36719_comb;
  wire [26:0] p8_add_36721_comb;
  wire [26:0] p8_add_36723_comb;
  wire [26:0] p8_add_36725_comb;
  wire [28:0] p8_concat_36743_comb;
  wire [18:0] p8_add_36727_comb;
  wire [4:0] p8_bit_slice_36728_comb;
  wire [28:0] p8_concat_36744_comb;
  wire [18:0] p8_add_36730_comb;
  wire [4:0] p8_bit_slice_36731_comb;
  wire [28:0] p8_concat_36745_comb;
  wire [18:0] p8_add_36733_comb;
  wire [4:0] p8_bit_slice_36734_comb;
  wire [28:0] p8_concat_36746_comb;
  wire [18:0] p8_add_36736_comb;
  wire [4:0] p8_bit_slice_36737_comb;
  wire [31:0] p8_sign_ext_36755_comb;
  wire [23:0] p8_bit_slice_36729_comb;
  wire [31:0] p8_sign_ext_36757_comb;
  wire [23:0] p8_bit_slice_36732_comb;
  wire [31:0] p8_sign_ext_36759_comb;
  wire [23:0] p8_bit_slice_36735_comb;
  wire [31:0] p8_sign_ext_36761_comb;
  wire [23:0] p8_bit_slice_36738_comb;
  wire [18:0] p8_add_36763_comb;
  wire [18:0] p8_add_36765_comb;
  wire [18:0] p8_add_36767_comb;
  wire [18:0] p8_add_36769_comb;
  wire [23:0] p8_add_36772_comb;
  wire [23:0] p8_add_36774_comb;
  wire [23:0] p8_add_36776_comb;
  wire [23:0] p8_add_36778_comb;
  wire [23:0] p8_bit_slice_36779_comb;
  wire [23:0] p8_bit_slice_36780_comb;
  wire [23:0] p8_bit_slice_36781_comb;
  wire [23:0] p8_bit_slice_36782_comb;
  wire [23:0] p8_add_36791_comb;
  wire [23:0] p8_add_36793_comb;
  wire [23:0] p8_add_36795_comb;
  wire [23:0] p8_add_36797_comb;
  wire [23:0] p8_add_36803_comb;
  wire [23:0] p8_add_36805_comb;
  wire [23:0] p8_add_36807_comb;
  wire [23:0] p8_add_36809_comb;
  wire [31:0] p8_concat_36811_comb;
  wire [31:0] p8_concat_36812_comb;
  wire [31:0] p8_concat_36813_comb;
  wire [31:0] p8_concat_36814_comb;
  wire [31:0] p8_sub_36815_comb;
  wire [31:0] p8_sub_36816_comb;
  wire [31:0] p8_sub_36817_comb;
  wire [31:0] p8_sub_36818_comb;
  wire [31:0] p8_add_36820_comb;
  wire [31:0] p8_add_36822_comb;
  wire [31:0] p8_add_36824_comb;
  wire [31:0] p8_add_36826_comb;
  wire [31:0] p8_umul_36659_comb;
  wire [31:0] p8_umul_36660_comb;
  wire [31:0] p8_umul_36661_comb;
  wire [31:0] p8_umul_36662_comb;
  wire [31:0] p8_umul_36692_comb;
  wire [31:0] p8_umul_36694_comb;
  wire [31:0] p8_umul_36696_comb;
  wire [31:0] p8_umul_36698_comb;
  wire [31:0] p8_add_36827_comb;
  wire [31:0] p8_add_36828_comb;
  wire [31:0] p8_add_36829_comb;
  wire [31:0] p8_add_36830_comb;
  wire [31:0] p8_add_36831_comb;
  wire [31:0] p8_add_36832_comb;
  wire [31:0] p8_add_36833_comb;
  wire [31:0] p8_add_36834_comb;
  wire [31:0] p8_sub_36835_comb;
  wire [31:0] p8_sub_36836_comb;
  wire [31:0] p8_sub_36837_comb;
  wire [31:0] p8_sub_36838_comb;
  wire [31:0] p8_sub_36839_comb;
  wire [31:0] p8_sub_36840_comb;
  wire [31:0] p8_sub_36841_comb;
  wire [31:0] p8_sub_36842_comb;
  wire [31:0] p8_sub_36691_comb;
  wire [31:0] p8_sub_36693_comb;
  wire [31:0] p8_sub_36695_comb;
  wire [31:0] p8_sub_36697_comb;
  wire [17:0] p8_bit_slice_36843_comb;
  wire [17:0] p8_bit_slice_36844_comb;
  wire [17:0] p8_bit_slice_36845_comb;
  wire [17:0] p8_bit_slice_36846_comb;
  wire [17:0] p8_bit_slice_36847_comb;
  wire [17:0] p8_bit_slice_36848_comb;
  wire [17:0] p8_bit_slice_36849_comb;
  wire [17:0] p8_bit_slice_36850_comb;
  wire [17:0] p8_bit_slice_36851_comb;
  wire [17:0] p8_bit_slice_36852_comb;
  wire [17:0] p8_bit_slice_36853_comb;
  wire [17:0] p8_bit_slice_36854_comb;
  wire [17:0] p8_bit_slice_36855_comb;
  wire [17:0] p8_bit_slice_36856_comb;
  wire [17:0] p8_bit_slice_36857_comb;
  wire [17:0] p8_bit_slice_36858_comb;
  wire [24:0] p8_add_36687_comb;
  wire [24:0] p8_add_36688_comb;
  wire [24:0] p8_add_36689_comb;
  wire [24:0] p8_add_36690_comb;
  wire [24:0] p8_add_36739_comb;
  wire [24:0] p8_add_36740_comb;
  wire [24:0] p8_add_36741_comb;
  wire [24:0] p8_add_36742_comb;
  assign p8_add_36663_comb = p7_bit_slice_36199 + 30'h0000_0001;
  assign p8_add_36665_comb = p7_bit_slice_36200 + 30'h0000_0001;
  assign p8_add_36667_comb = p7_bit_slice_36201 + 30'h0000_0001;
  assign p8_add_36669_comb = p7_bit_slice_36202 + 30'h0000_0001;
  assign p8_add_36719_comb = p7_bit_slice_36299 + p8_add_36663_comb[29:3];
  assign p8_add_36721_comb = p7_bit_slice_36300 + p8_add_36665_comb[29:3];
  assign p8_add_36723_comb = p7_bit_slice_36301 + p8_add_36667_comb[29:3];
  assign p8_add_36725_comb = p7_bit_slice_36302 + p8_add_36669_comb[29:3];
  assign p8_concat_36743_comb = {p8_add_36719_comb, p8_add_36663_comb[2:1]};
  assign p8_add_36727_comb = p7_sub_36287[31:13] + 19'h0_0001;
  assign p8_bit_slice_36728_comb = p7_sub_36287[12:8];
  assign p8_concat_36744_comb = {p8_add_36721_comb, p8_add_36665_comb[2:1]};
  assign p8_add_36730_comb = p7_sub_36290[31:13] + 19'h0_0001;
  assign p8_bit_slice_36731_comb = p7_sub_36290[12:8];
  assign p8_concat_36745_comb = {p8_add_36723_comb, p8_add_36667_comb[2:1]};
  assign p8_add_36733_comb = p7_sub_36293[31:13] + 19'h0_0001;
  assign p8_bit_slice_36734_comb = p7_sub_36293[12:8];
  assign p8_concat_36746_comb = {p8_add_36725_comb, p8_add_36669_comb[2:1]};
  assign p8_add_36736_comb = p7_sub_36296[31:13] + 19'h0_0001;
  assign p8_bit_slice_36737_comb = p7_sub_36296[12:8];
  assign p8_sign_ext_36755_comb = {{3{p8_concat_36743_comb[28]}}, p8_concat_36743_comb};
  assign p8_bit_slice_36729_comb = p7_sub_36303[31:8];
  assign p8_sign_ext_36757_comb = {{3{p8_concat_36744_comb[28]}}, p8_concat_36744_comb};
  assign p8_bit_slice_36732_comb = p7_sub_36304[31:8];
  assign p8_sign_ext_36759_comb = {{3{p8_concat_36745_comb[28]}}, p8_concat_36745_comb};
  assign p8_bit_slice_36735_comb = p7_sub_36305[31:8];
  assign p8_sign_ext_36761_comb = {{3{p8_concat_36746_comb[28]}}, p8_concat_36746_comb};
  assign p8_bit_slice_36738_comb = p7_sub_36306[31:8];
  assign p8_add_36763_comb = p7_sub_36303[31:13] + 19'h0_0001;
  assign p8_add_36765_comb = p7_sub_36304[31:13] + 19'h0_0001;
  assign p8_add_36767_comb = p7_sub_36305[31:13] + 19'h0_0001;
  assign p8_add_36769_comb = p7_sub_36306[31:13] + 19'h0_0001;
  assign p8_add_36772_comb = p8_bit_slice_36729_comb + {p8_add_36727_comb, p8_bit_slice_36728_comb};
  assign p8_add_36774_comb = p8_bit_slice_36732_comb + {p8_add_36730_comb, p8_bit_slice_36731_comb};
  assign p8_add_36776_comb = p8_bit_slice_36735_comb + {p8_add_36733_comb, p8_bit_slice_36734_comb};
  assign p8_add_36778_comb = p8_bit_slice_36738_comb + {p8_add_36736_comb, p8_bit_slice_36737_comb};
  assign p8_bit_slice_36779_comb = p7_sub_36287[31:8];
  assign p8_bit_slice_36780_comb = p7_sub_36290[31:8];
  assign p8_bit_slice_36781_comb = p7_sub_36293[31:8];
  assign p8_bit_slice_36782_comb = p7_sub_36296[31:8];
  assign p8_add_36791_comb = p8_sign_ext_36755_comb[31:8] + p8_add_36772_comb;
  assign p8_add_36793_comb = p8_sign_ext_36757_comb[31:8] + p8_add_36774_comb;
  assign p8_add_36795_comb = p8_sign_ext_36759_comb[31:8] + p8_add_36776_comb;
  assign p8_add_36797_comb = p8_sign_ext_36761_comb[31:8] + p8_add_36778_comb;
  assign p8_add_36803_comb = {p8_add_36763_comb, p7_sub_36303[12:8]} + p8_bit_slice_36779_comb;
  assign p8_add_36805_comb = {p8_add_36765_comb, p7_sub_36304[12:8]} + p8_bit_slice_36780_comb;
  assign p8_add_36807_comb = {p8_add_36767_comb, p7_sub_36305[12:8]} + p8_bit_slice_36781_comb;
  assign p8_add_36809_comb = {p8_add_36769_comb, p7_sub_36306[12:8]} + p8_bit_slice_36782_comb;
  assign p8_concat_36811_comb = {p8_add_36791_comb, p8_add_36719_comb[5:0], p8_add_36663_comb[2:1]};
  assign p8_concat_36812_comb = {p8_add_36793_comb, p8_add_36721_comb[5:0], p8_add_36665_comb[2:1]};
  assign p8_concat_36813_comb = {p8_add_36795_comb, p8_add_36723_comb[5:0], p8_add_36667_comb[2:1]};
  assign p8_concat_36814_comb = {p8_add_36797_comb, p8_add_36725_comb[5:0], p8_add_36669_comb[2:1]};
  assign p8_sub_36815_comb = {p8_add_36772_comb, 8'h00} - p8_sign_ext_36755_comb;
  assign p8_sub_36816_comb = {p8_add_36774_comb, 8'h00} - p8_sign_ext_36757_comb;
  assign p8_sub_36817_comb = {p8_add_36776_comb, 8'h00} - p8_sign_ext_36759_comb;
  assign p8_sub_36818_comb = {p8_add_36778_comb, 8'h00} - p8_sign_ext_36761_comb;
  assign p8_add_36820_comb = p8_sign_ext_36755_comb + p7_add_36431;
  assign p8_add_36822_comb = p8_sign_ext_36757_comb + p7_add_36432;
  assign p8_add_36824_comb = p8_sign_ext_36759_comb + p7_add_36433;
  assign p8_add_36826_comb = p8_sign_ext_36761_comb + p7_add_36434;
  assign p8_umul_36659_comb = umul32b_32b_x_8b(p7_sub_36195, 8'hb5);
  assign p8_umul_36660_comb = umul32b_32b_x_8b(p7_sub_36196, 8'hb5);
  assign p8_umul_36661_comb = umul32b_32b_x_8b(p7_sub_36197, 8'hb5);
  assign p8_umul_36662_comb = umul32b_32b_x_8b(p7_sub_36198, 8'hb5);
  assign p8_umul_36692_comb = umul32b_32b_x_8b(p7_sub_36276, 8'hb5);
  assign p8_umul_36694_comb = umul32b_32b_x_8b(p7_sub_36278, 8'hb5);
  assign p8_umul_36696_comb = umul32b_32b_x_8b(p7_sub_36280, 8'hb5);
  assign p8_umul_36698_comb = umul32b_32b_x_8b(p7_sub_36282, 8'hb5);
  assign p8_add_36827_comb = p7_add_36455 + p8_concat_36811_comb;
  assign p8_add_36828_comb = p7_add_36456 + p8_concat_36812_comb;
  assign p8_add_36829_comb = p7_add_36457 + p8_concat_36813_comb;
  assign p8_add_36830_comb = p7_add_36458 + p8_concat_36814_comb;
  assign p8_add_36831_comb = p8_sub_36815_comb + p7_add_36431;
  assign p8_add_36832_comb = p8_sub_36816_comb + p7_add_36432;
  assign p8_add_36833_comb = p8_sub_36817_comb + p7_add_36433;
  assign p8_add_36834_comb = p8_sub_36818_comb + p7_add_36434;
  assign p8_sub_36835_comb = {p8_add_36803_comb, 8'h00} - p8_add_36820_comb;
  assign p8_sub_36836_comb = {p8_add_36805_comb, 8'h00} - p8_add_36822_comb;
  assign p8_sub_36837_comb = {p8_add_36807_comb, 8'h00} - p8_add_36824_comb;
  assign p8_sub_36838_comb = {p8_add_36809_comb, 8'h00} - p8_add_36826_comb;
  assign p8_sub_36839_comb = p8_concat_36811_comb - p7_add_36455;
  assign p8_sub_36840_comb = p8_concat_36812_comb - p7_add_36456;
  assign p8_sub_36841_comb = p8_concat_36813_comb - p7_add_36457;
  assign p8_sub_36842_comb = p8_concat_36814_comb - p7_add_36458;
  assign p8_sub_36691_comb = {p8_add_36663_comb, 2'h0} - p7_umul_36275;
  assign p8_sub_36693_comb = {p8_add_36665_comb, 2'h0} - p7_umul_36277;
  assign p8_sub_36695_comb = {p8_add_36667_comb, 2'h0} - p7_umul_36279;
  assign p8_sub_36697_comb = {p8_add_36669_comb, 2'h0} - p7_umul_36281;
  assign p8_bit_slice_36843_comb = p8_add_36827_comb[31:14];
  assign p8_bit_slice_36844_comb = p8_add_36828_comb[31:14];
  assign p8_bit_slice_36845_comb = p8_add_36829_comb[31:14];
  assign p8_bit_slice_36846_comb = p8_add_36830_comb[31:14];
  assign p8_bit_slice_36847_comb = p8_add_36831_comb[31:14];
  assign p8_bit_slice_36848_comb = p8_add_36832_comb[31:14];
  assign p8_bit_slice_36849_comb = p8_add_36833_comb[31:14];
  assign p8_bit_slice_36850_comb = p8_add_36834_comb[31:14];
  assign p8_bit_slice_36851_comb = p8_sub_36835_comb[31:14];
  assign p8_bit_slice_36852_comb = p8_sub_36836_comb[31:14];
  assign p8_bit_slice_36853_comb = p8_sub_36837_comb[31:14];
  assign p8_bit_slice_36854_comb = p8_sub_36838_comb[31:14];
  assign p8_bit_slice_36855_comb = p8_sub_36839_comb[31:14];
  assign p8_bit_slice_36856_comb = p8_sub_36840_comb[31:14];
  assign p8_bit_slice_36857_comb = p8_sub_36841_comb[31:14];
  assign p8_bit_slice_36858_comb = p8_sub_36842_comb[31:14];
  assign p8_add_36687_comb = p8_umul_36659_comb[31:7] + 25'h000_0001;
  assign p8_add_36688_comb = p8_umul_36660_comb[31:7] + 25'h000_0001;
  assign p8_add_36689_comb = p8_umul_36661_comb[31:7] + 25'h000_0001;
  assign p8_add_36690_comb = p8_umul_36662_comb[31:7] + 25'h000_0001;
  assign p8_add_36739_comb = p8_umul_36692_comb[31:7] + 25'h000_0001;
  assign p8_add_36740_comb = p8_umul_36694_comb[31:7] + 25'h000_0001;
  assign p8_add_36741_comb = p8_umul_36696_comb[31:7] + 25'h000_0001;
  assign p8_add_36742_comb = p8_umul_36698_comb[31:7] + 25'h000_0001;

  // Registers for pipe stage 8:
  reg [31:0] p8_sub_36691;
  reg [31:0] p8_sub_36693;
  reg [31:0] p8_sub_36695;
  reg [31:0] p8_sub_36697;
  reg [4:0] p8_bit_slice_36728;
  reg [23:0] p8_bit_slice_36729;
  reg [4:0] p8_bit_slice_36731;
  reg [23:0] p8_bit_slice_36732;
  reg [4:0] p8_bit_slice_36734;
  reg [23:0] p8_bit_slice_36735;
  reg [4:0] p8_bit_slice_36737;
  reg [23:0] p8_bit_slice_36738;
  reg [23:0] p8_bit_slice_36779;
  reg [23:0] p8_bit_slice_36780;
  reg [23:0] p8_bit_slice_36781;
  reg [23:0] p8_bit_slice_36782;
  reg [17:0] p8_bit_slice_35831;
  reg [17:0] p8_bit_slice_36843;
  reg [17:0] p8_bit_slice_36844;
  reg [17:0] p8_bit_slice_35832;
  reg [17:0] p8_bit_slice_35833;
  reg [17:0] p8_bit_slice_36845;
  reg [17:0] p8_bit_slice_36846;
  reg [17:0] p8_bit_slice_35834;
  reg [17:0] p8_bit_slice_36499;
  reg [17:0] p8_bit_slice_36500;
  reg [17:0] p8_bit_slice_36501;
  reg [17:0] p8_bit_slice_36502;
  reg [17:0] p8_bit_slice_36503;
  reg [17:0] p8_bit_slice_36504;
  reg [17:0] p8_bit_slice_36505;
  reg [17:0] p8_bit_slice_36506;
  reg [17:0] p8_bit_slice_35835;
  reg [17:0] p8_bit_slice_36847;
  reg [17:0] p8_bit_slice_36848;
  reg [17:0] p8_bit_slice_35836;
  reg [17:0] p8_bit_slice_35837;
  reg [17:0] p8_bit_slice_36849;
  reg [17:0] p8_bit_slice_36850;
  reg [17:0] p8_bit_slice_35838;
  reg [17:0] p8_bit_slice_35839;
  reg [17:0] p8_bit_slice_36851;
  reg [17:0] p8_bit_slice_36852;
  reg [17:0] p8_bit_slice_35840;
  reg [17:0] p8_bit_slice_35841;
  reg [17:0] p8_bit_slice_36853;
  reg [17:0] p8_bit_slice_36854;
  reg [17:0] p8_bit_slice_35842;
  reg [17:0] p8_bit_slice_36507;
  reg [17:0] p8_bit_slice_36508;
  reg [17:0] p8_bit_slice_36509;
  reg [17:0] p8_bit_slice_36510;
  reg [17:0] p8_bit_slice_36511;
  reg [17:0] p8_bit_slice_36512;
  reg [17:0] p8_bit_slice_36513;
  reg [17:0] p8_bit_slice_36514;
  reg [17:0] p8_bit_slice_35843;
  reg [17:0] p8_bit_slice_36855;
  reg [17:0] p8_bit_slice_36856;
  reg [17:0] p8_bit_slice_35844;
  reg [17:0] p8_bit_slice_35845;
  reg [17:0] p8_bit_slice_36857;
  reg [17:0] p8_bit_slice_36858;
  reg [17:0] p8_bit_slice_35846;
  reg [24:0] p8_add_36687;
  reg [24:0] p8_add_36688;
  reg [24:0] p8_add_36689;
  reg [24:0] p8_add_36690;
  reg [18:0] p8_add_36727;
  reg [18:0] p8_add_36730;
  reg [18:0] p8_add_36733;
  reg [18:0] p8_add_36736;
  reg [24:0] p8_add_36739;
  reg [24:0] p8_add_36740;
  reg [24:0] p8_add_36741;
  reg [24:0] p8_add_36742;
  always_ff @ (posedge clk) begin
    p8_sub_36691 <= p8_sub_36691_comb;
    p8_sub_36693 <= p8_sub_36693_comb;
    p8_sub_36695 <= p8_sub_36695_comb;
    p8_sub_36697 <= p8_sub_36697_comb;
    p8_bit_slice_36728 <= p8_bit_slice_36728_comb;
    p8_bit_slice_36729 <= p8_bit_slice_36729_comb;
    p8_bit_slice_36731 <= p8_bit_slice_36731_comb;
    p8_bit_slice_36732 <= p8_bit_slice_36732_comb;
    p8_bit_slice_36734 <= p8_bit_slice_36734_comb;
    p8_bit_slice_36735 <= p8_bit_slice_36735_comb;
    p8_bit_slice_36737 <= p8_bit_slice_36737_comb;
    p8_bit_slice_36738 <= p8_bit_slice_36738_comb;
    p8_bit_slice_36779 <= p8_bit_slice_36779_comb;
    p8_bit_slice_36780 <= p8_bit_slice_36780_comb;
    p8_bit_slice_36781 <= p8_bit_slice_36781_comb;
    p8_bit_slice_36782 <= p8_bit_slice_36782_comb;
    p8_bit_slice_35831 <= p7_bit_slice_35831;
    p8_bit_slice_36843 <= p8_bit_slice_36843_comb;
    p8_bit_slice_36844 <= p8_bit_slice_36844_comb;
    p8_bit_slice_35832 <= p7_bit_slice_35832;
    p8_bit_slice_35833 <= p7_bit_slice_35833;
    p8_bit_slice_36845 <= p8_bit_slice_36845_comb;
    p8_bit_slice_36846 <= p8_bit_slice_36846_comb;
    p8_bit_slice_35834 <= p7_bit_slice_35834;
    p8_bit_slice_36499 <= p7_bit_slice_36499;
    p8_bit_slice_36500 <= p7_bit_slice_36500;
    p8_bit_slice_36501 <= p7_bit_slice_36501;
    p8_bit_slice_36502 <= p7_bit_slice_36502;
    p8_bit_slice_36503 <= p7_bit_slice_36503;
    p8_bit_slice_36504 <= p7_bit_slice_36504;
    p8_bit_slice_36505 <= p7_bit_slice_36505;
    p8_bit_slice_36506 <= p7_bit_slice_36506;
    p8_bit_slice_35835 <= p7_bit_slice_35835;
    p8_bit_slice_36847 <= p8_bit_slice_36847_comb;
    p8_bit_slice_36848 <= p8_bit_slice_36848_comb;
    p8_bit_slice_35836 <= p7_bit_slice_35836;
    p8_bit_slice_35837 <= p7_bit_slice_35837;
    p8_bit_slice_36849 <= p8_bit_slice_36849_comb;
    p8_bit_slice_36850 <= p8_bit_slice_36850_comb;
    p8_bit_slice_35838 <= p7_bit_slice_35838;
    p8_bit_slice_35839 <= p7_bit_slice_35839;
    p8_bit_slice_36851 <= p8_bit_slice_36851_comb;
    p8_bit_slice_36852 <= p8_bit_slice_36852_comb;
    p8_bit_slice_35840 <= p7_bit_slice_35840;
    p8_bit_slice_35841 <= p7_bit_slice_35841;
    p8_bit_slice_36853 <= p8_bit_slice_36853_comb;
    p8_bit_slice_36854 <= p8_bit_slice_36854_comb;
    p8_bit_slice_35842 <= p7_bit_slice_35842;
    p8_bit_slice_36507 <= p7_bit_slice_36507;
    p8_bit_slice_36508 <= p7_bit_slice_36508;
    p8_bit_slice_36509 <= p7_bit_slice_36509;
    p8_bit_slice_36510 <= p7_bit_slice_36510;
    p8_bit_slice_36511 <= p7_bit_slice_36511;
    p8_bit_slice_36512 <= p7_bit_slice_36512;
    p8_bit_slice_36513 <= p7_bit_slice_36513;
    p8_bit_slice_36514 <= p7_bit_slice_36514;
    p8_bit_slice_35843 <= p7_bit_slice_35843;
    p8_bit_slice_36855 <= p8_bit_slice_36855_comb;
    p8_bit_slice_36856 <= p8_bit_slice_36856_comb;
    p8_bit_slice_35844 <= p7_bit_slice_35844;
    p8_bit_slice_35845 <= p7_bit_slice_35845;
    p8_bit_slice_36857 <= p8_bit_slice_36857_comb;
    p8_bit_slice_36858 <= p8_bit_slice_36858_comb;
    p8_bit_slice_35846 <= p7_bit_slice_35846;
    p8_add_36687 <= p8_add_36687_comb;
    p8_add_36688 <= p8_add_36688_comb;
    p8_add_36689 <= p8_add_36689_comb;
    p8_add_36690 <= p8_add_36690_comb;
    p8_add_36727 <= p8_add_36727_comb;
    p8_add_36730 <= p8_add_36730_comb;
    p8_add_36733 <= p8_add_36733_comb;
    p8_add_36736 <= p8_add_36736_comb;
    p8_add_36739 <= p8_add_36739_comb;
    p8_add_36740 <= p8_add_36740_comb;
    p8_add_36741 <= p8_add_36741_comb;
    p8_add_36742 <= p8_add_36742_comb;
  end

  // ===== Pipe stage 9:
  wire [23:0] p9_bit_slice_37011_comb;
  wire [23:0] p9_bit_slice_37012_comb;
  wire [23:0] p9_bit_slice_37013_comb;
  wire [23:0] p9_bit_slice_37014_comb;
  wire [28:0] p9_bit_slice_37015_comb;
  wire [28:0] p9_bit_slice_37016_comb;
  wire [28:0] p9_bit_slice_37017_comb;
  wire [28:0] p9_bit_slice_37018_comb;
  wire [31:0] p9_sign_ext_37027_comb;
  wire [31:0] p9_sign_ext_37028_comb;
  wire [31:0] p9_sign_ext_37029_comb;
  wire [31:0] p9_sign_ext_37030_comb;
  wire [31:0] p9_sign_ext_37031_comb;
  wire [31:0] p9_sign_ext_37032_comb;
  wire [31:0] p9_sign_ext_37033_comb;
  wire [31:0] p9_sign_ext_37034_comb;
  wire [31:0] p9_concat_37035_comb;
  wire [31:0] p9_concat_37037_comb;
  wire [31:0] p9_concat_37039_comb;
  wire [31:0] p9_concat_37041_comb;
  wire [23:0] p9_bit_slice_37053_comb;
  wire [23:0] p9_bit_slice_37056_comb;
  wire [23:0] p9_bit_slice_37059_comb;
  wire [23:0] p9_bit_slice_37062_comb;
  wire [31:0] p9_sub_37063_comb;
  wire [31:0] p9_sub_37064_comb;
  wire [31:0] p9_sub_37065_comb;
  wire [31:0] p9_sub_37066_comb;
  wire [18:0] p9_add_37067_comb;
  wire [18:0] p9_add_37069_comb;
  wire [18:0] p9_add_37071_comb;
  wire [18:0] p9_add_37073_comb;
  wire [31:0] p9_add_37075_comb;
  wire [31:0] p9_add_37076_comb;
  wire [31:0] p9_add_37077_comb;
  wire [31:0] p9_add_37078_comb;
  wire [18:0] p9_add_37079_comb;
  wire [31:0] p9_sign_ext_37081_comb;
  wire [18:0] p9_add_37082_comb;
  wire [31:0] p9_sign_ext_37084_comb;
  wire [18:0] p9_add_37085_comb;
  wire [31:0] p9_sign_ext_37087_comb;
  wire [18:0] p9_add_37088_comb;
  wire [31:0] p9_sign_ext_37090_comb;
  wire [23:0] p9_add_37115_comb;
  wire [23:0] p9_add_37117_comb;
  wire [23:0] p9_add_37119_comb;
  wire [23:0] p9_add_37121_comb;
  wire [23:0] p9_add_37123_comb;
  wire [23:0] p9_add_37125_comb;
  wire [23:0] p9_add_37126_comb;
  wire [23:0] p9_add_37128_comb;
  wire [23:0] p9_add_37129_comb;
  wire [23:0] p9_add_37131_comb;
  wire [23:0] p9_add_37132_comb;
  wire [23:0] p9_add_37134_comb;
  wire [23:0] p9_add_37135_comb;
  wire [23:0] p9_add_37137_comb;
  wire [23:0] p9_add_37139_comb;
  wire [23:0] p9_add_37141_comb;
  wire [23:0] p9_add_37143_comb;
  wire [23:0] p9_add_37144_comb;
  wire [23:0] p9_add_37146_comb;
  wire [23:0] p9_add_37147_comb;
  wire [23:0] p9_add_37149_comb;
  wire [23:0] p9_add_37150_comb;
  wire [23:0] p9_add_37152_comb;
  wire [23:0] p9_add_37153_comb;
  wire [31:0] p9_add_37179_comb;
  wire [31:0] p9_add_37180_comb;
  wire [31:0] p9_add_37181_comb;
  wire [31:0] p9_add_37182_comb;
  wire [31:0] p9_sub_37183_comb;
  wire [31:0] p9_sub_37184_comb;
  wire [31:0] p9_sub_37185_comb;
  wire [31:0] p9_sub_37186_comb;
  wire [31:0] p9_sub_37187_comb;
  wire [31:0] p9_sub_37188_comb;
  wire [31:0] p9_sub_37189_comb;
  wire [31:0] p9_sub_37190_comb;
  wire [31:0] p9_sub_37191_comb;
  wire [31:0] p9_sub_37192_comb;
  wire [31:0] p9_sub_37193_comb;
  wire [31:0] p9_sub_37194_comb;
  wire [17:0] p9_bit_slice_37195_comb;
  wire [17:0] p9_bit_slice_37196_comb;
  wire [17:0] p9_bit_slice_37197_comb;
  wire [17:0] p9_bit_slice_37198_comb;
  wire [17:0] p9_bit_slice_37199_comb;
  wire [17:0] p9_bit_slice_37200_comb;
  wire [17:0] p9_bit_slice_37201_comb;
  wire [17:0] p9_bit_slice_37202_comb;
  wire [17:0] p9_bit_slice_37203_comb;
  wire [17:0] p9_bit_slice_37204_comb;
  wire [17:0] p9_bit_slice_37205_comb;
  wire [17:0] p9_bit_slice_37206_comb;
  wire [17:0] p9_bit_slice_37207_comb;
  wire [17:0] p9_bit_slice_37208_comb;
  wire [17:0] p9_bit_slice_37209_comb;
  wire [17:0] p9_bit_slice_37210_comb;
  wire [31:0] p9_array_37275_comb[64];
  assign p9_bit_slice_37011_comb = p8_add_36687[24:1];
  assign p9_bit_slice_37012_comb = p8_add_36688[24:1];
  assign p9_bit_slice_37013_comb = p8_add_36689[24:1];
  assign p9_bit_slice_37014_comb = p8_add_36690[24:1];
  assign p9_bit_slice_37015_comb = p8_sub_36691[31:3];
  assign p9_bit_slice_37016_comb = p8_sub_36693[31:3];
  assign p9_bit_slice_37017_comb = p8_sub_36695[31:3];
  assign p9_bit_slice_37018_comb = p8_sub_36697[31:3];
  assign p9_sign_ext_37027_comb = {{8{p9_bit_slice_37011_comb[23]}}, p9_bit_slice_37011_comb};
  assign p9_sign_ext_37028_comb = {{8{p9_bit_slice_37012_comb[23]}}, p9_bit_slice_37012_comb};
  assign p9_sign_ext_37029_comb = {{8{p9_bit_slice_37013_comb[23]}}, p9_bit_slice_37013_comb};
  assign p9_sign_ext_37030_comb = {{8{p9_bit_slice_37014_comb[23]}}, p9_bit_slice_37014_comb};
  assign p9_sign_ext_37031_comb = {{3{p9_bit_slice_37015_comb[28]}}, p9_bit_slice_37015_comb};
  assign p9_sign_ext_37032_comb = {{3{p9_bit_slice_37016_comb[28]}}, p9_bit_slice_37016_comb};
  assign p9_sign_ext_37033_comb = {{3{p9_bit_slice_37017_comb[28]}}, p9_bit_slice_37017_comb};
  assign p9_sign_ext_37034_comb = {{3{p9_bit_slice_37018_comb[28]}}, p9_bit_slice_37018_comb};
  assign p9_concat_37035_comb = {p8_add_36727, p8_bit_slice_36728, 8'h00};
  assign p9_concat_37037_comb = {p8_add_36730, p8_bit_slice_36731, 8'h00};
  assign p9_concat_37039_comb = {p8_add_36733, p8_bit_slice_36734, 8'h00};
  assign p9_concat_37041_comb = {p8_add_36736, p8_bit_slice_36737, 8'h00};
  assign p9_bit_slice_37053_comb = p8_add_36739[24:1];
  assign p9_bit_slice_37056_comb = p8_add_36740[24:1];
  assign p9_bit_slice_37059_comb = p8_add_36741[24:1];
  assign p9_bit_slice_37062_comb = p8_add_36742[24:1];
  assign p9_sub_37063_comb = p9_concat_37035_comb - {p8_bit_slice_36729, 8'h00};
  assign p9_sub_37064_comb = p9_concat_37037_comb - {p8_bit_slice_36732, 8'h00};
  assign p9_sub_37065_comb = p9_concat_37039_comb - {p8_bit_slice_36735, 8'h00};
  assign p9_sub_37066_comb = p9_concat_37041_comb - {p8_bit_slice_36738, 8'h00};
  assign p9_add_37067_comb = p9_sign_ext_37027_comb[31:13] + 19'h0_0001;
  assign p9_add_37069_comb = p9_sign_ext_37028_comb[31:13] + 19'h0_0001;
  assign p9_add_37071_comb = p9_sign_ext_37029_comb[31:13] + 19'h0_0001;
  assign p9_add_37073_comb = p9_sign_ext_37030_comb[31:13] + 19'h0_0001;
  assign p9_add_37075_comb = p9_sign_ext_37027_comb + p9_sign_ext_37031_comb;
  assign p9_add_37076_comb = p9_sign_ext_37028_comb + p9_sign_ext_37032_comb;
  assign p9_add_37077_comb = p9_sign_ext_37029_comb + p9_sign_ext_37033_comb;
  assign p9_add_37078_comb = p9_sign_ext_37030_comb + p9_sign_ext_37034_comb;
  assign p9_add_37079_comb = p9_sign_ext_37031_comb[31:13] + 19'h0_0001;
  assign p9_sign_ext_37081_comb = {{8{p9_bit_slice_37053_comb[23]}}, p9_bit_slice_37053_comb};
  assign p9_add_37082_comb = p9_sign_ext_37032_comb[31:13] + 19'h0_0001;
  assign p9_sign_ext_37084_comb = {{8{p9_bit_slice_37056_comb[23]}}, p9_bit_slice_37056_comb};
  assign p9_add_37085_comb = p9_sign_ext_37033_comb[31:13] + 19'h0_0001;
  assign p9_sign_ext_37087_comb = {{8{p9_bit_slice_37059_comb[23]}}, p9_bit_slice_37059_comb};
  assign p9_add_37088_comb = p9_sign_ext_37034_comb[31:13] + 19'h0_0001;
  assign p9_sign_ext_37090_comb = {{8{p9_bit_slice_37062_comb[23]}}, p9_bit_slice_37062_comb};
  assign p9_add_37115_comb = p9_sign_ext_37031_comb[31:8] + p9_sub_37063_comb[31:8];
  assign p9_add_37117_comb = p9_sign_ext_37032_comb[31:8] + p9_sub_37064_comb[31:8];
  assign p9_add_37119_comb = p9_sign_ext_37033_comb[31:8] + p9_sub_37065_comb[31:8];
  assign p9_add_37121_comb = p9_sign_ext_37034_comb[31:8] + p9_sub_37066_comb[31:8];
  assign p9_add_37123_comb = {p9_add_37067_comb, p8_add_36687[13:9]} + p8_bit_slice_36779;
  assign p9_add_37125_comb = p9_sign_ext_37031_comb[31:8] + p8_bit_slice_36729;
  assign p9_add_37126_comb = {p9_add_37069_comb, p8_add_36688[13:9]} + p8_bit_slice_36780;
  assign p9_add_37128_comb = p9_sign_ext_37032_comb[31:8] + p8_bit_slice_36732;
  assign p9_add_37129_comb = {p9_add_37071_comb, p8_add_36689[13:9]} + p8_bit_slice_36781;
  assign p9_add_37131_comb = p9_sign_ext_37033_comb[31:8] + p8_bit_slice_36735;
  assign p9_add_37132_comb = {p9_add_37073_comb, p8_add_36690[13:9]} + p8_bit_slice_36782;
  assign p9_add_37134_comb = p9_sign_ext_37034_comb[31:8] + p8_bit_slice_36738;
  assign p9_add_37135_comb = p9_add_37075_comb[31:8] + p8_bit_slice_36729;
  assign p9_add_37137_comb = p9_add_37076_comb[31:8] + p8_bit_slice_36732;
  assign p9_add_37139_comb = p9_add_37077_comb[31:8] + p8_bit_slice_36735;
  assign p9_add_37141_comb = p9_add_37078_comb[31:8] + p8_bit_slice_36738;
  assign p9_add_37143_comb = {p9_add_37079_comb, p8_sub_36691[15:11]} + p8_bit_slice_36779;
  assign p9_add_37144_comb = p9_sign_ext_37081_comb[31:8] + p8_bit_slice_36729;
  assign p9_add_37146_comb = {p9_add_37082_comb, p8_sub_36693[15:11]} + p8_bit_slice_36780;
  assign p9_add_37147_comb = p9_sign_ext_37084_comb[31:8] + p8_bit_slice_36732;
  assign p9_add_37149_comb = {p9_add_37085_comb, p8_sub_36695[15:11]} + p8_bit_slice_36781;
  assign p9_add_37150_comb = p9_sign_ext_37087_comb[31:8] + p8_bit_slice_36735;
  assign p9_add_37152_comb = {p9_add_37088_comb, p8_sub_36697[15:11]} + p8_bit_slice_36782;
  assign p9_add_37153_comb = p9_sign_ext_37090_comb[31:8] + p8_bit_slice_36738;
  assign p9_add_37179_comb = p9_sign_ext_37081_comb + {p9_add_37115_comb, p8_sub_36691[10:3]};
  assign p9_add_37180_comb = p9_sign_ext_37084_comb + {p9_add_37117_comb, p8_sub_36693[10:3]};
  assign p9_add_37181_comb = p9_sign_ext_37087_comb + {p9_add_37119_comb, p8_sub_36695[10:3]};
  assign p9_add_37182_comb = p9_sign_ext_37090_comb + {p9_add_37121_comb, p8_sub_36697[10:3]};
  assign p9_sub_37183_comb = {p9_add_37123_comb, p8_add_36687[8:1]} - {p9_add_37125_comb, p8_sub_36691[10:3]};
  assign p9_sub_37184_comb = {p9_add_37126_comb, p8_add_36688[8:1]} - {p9_add_37128_comb, p8_sub_36693[10:3]};
  assign p9_sub_37185_comb = {p9_add_37129_comb, p8_add_36689[8:1]} - {p9_add_37131_comb, p8_sub_36695[10:3]};
  assign p9_sub_37186_comb = {p9_add_37132_comb, p8_add_36690[8:1]} - {p9_add_37134_comb, p8_sub_36697[10:3]};
  assign p9_sub_37187_comb = p9_concat_37035_comb - {p9_add_37135_comb, p9_add_37075_comb[7:0]};
  assign p9_sub_37188_comb = p9_concat_37037_comb - {p9_add_37137_comb, p9_add_37076_comb[7:0]};
  assign p9_sub_37189_comb = p9_concat_37039_comb - {p9_add_37139_comb, p9_add_37077_comb[7:0]};
  assign p9_sub_37190_comb = p9_concat_37041_comb - {p9_add_37141_comb, p9_add_37078_comb[7:0]};
  assign p9_sub_37191_comb = {p9_add_37143_comb, p8_sub_36691[10:3]} - {p9_add_37144_comb, p8_add_36739[8:1]};
  assign p9_sub_37192_comb = {p9_add_37146_comb, p8_sub_36693[10:3]} - {p9_add_37147_comb, p8_add_36740[8:1]};
  assign p9_sub_37193_comb = {p9_add_37149_comb, p8_sub_36695[10:3]} - {p9_add_37150_comb, p8_add_36741[8:1]};
  assign p9_sub_37194_comb = {p9_add_37152_comb, p8_sub_36697[10:3]} - {p9_add_37153_comb, p8_add_36742[8:1]};
  assign p9_bit_slice_37195_comb = p9_add_37179_comb[31:14];
  assign p9_bit_slice_37196_comb = p9_add_37180_comb[31:14];
  assign p9_bit_slice_37197_comb = p9_add_37181_comb[31:14];
  assign p9_bit_slice_37198_comb = p9_add_37182_comb[31:14];
  assign p9_bit_slice_37199_comb = p9_sub_37183_comb[31:14];
  assign p9_bit_slice_37200_comb = p9_sub_37184_comb[31:14];
  assign p9_bit_slice_37201_comb = p9_sub_37185_comb[31:14];
  assign p9_bit_slice_37202_comb = p9_sub_37186_comb[31:14];
  assign p9_bit_slice_37203_comb = p9_sub_37187_comb[31:14];
  assign p9_bit_slice_37204_comb = p9_sub_37188_comb[31:14];
  assign p9_bit_slice_37205_comb = p9_sub_37189_comb[31:14];
  assign p9_bit_slice_37206_comb = p9_sub_37190_comb[31:14];
  assign p9_bit_slice_37207_comb = p9_sub_37191_comb[31:14];
  assign p9_bit_slice_37208_comb = p9_sub_37192_comb[31:14];
  assign p9_bit_slice_37209_comb = p9_sub_37193_comb[31:14];
  assign p9_bit_slice_37210_comb = p9_sub_37194_comb[31:14];
  assign p9_array_37275_comb[0] = {{14{p8_bit_slice_35831[17]}}, p8_bit_slice_35831};
  assign p9_array_37275_comb[1] = {{14{p8_bit_slice_36843[17]}}, p8_bit_slice_36843};
  assign p9_array_37275_comb[2] = {{14{p8_bit_slice_36844[17]}}, p8_bit_slice_36844};
  assign p9_array_37275_comb[3] = {{14{p8_bit_slice_35832[17]}}, p8_bit_slice_35832};
  assign p9_array_37275_comb[4] = {{14{p8_bit_slice_35833[17]}}, p8_bit_slice_35833};
  assign p9_array_37275_comb[5] = {{14{p8_bit_slice_36845[17]}}, p8_bit_slice_36845};
  assign p9_array_37275_comb[6] = {{14{p8_bit_slice_36846[17]}}, p8_bit_slice_36846};
  assign p9_array_37275_comb[7] = {{14{p8_bit_slice_35834[17]}}, p8_bit_slice_35834};
  assign p9_array_37275_comb[8] = {{14{p8_bit_slice_36499[17]}}, p8_bit_slice_36499};
  assign p9_array_37275_comb[9] = {{14{p9_bit_slice_37195_comb[17]}}, p9_bit_slice_37195_comb};
  assign p9_array_37275_comb[10] = {{14{p9_bit_slice_37196_comb[17]}}, p9_bit_slice_37196_comb};
  assign p9_array_37275_comb[11] = {{14{p8_bit_slice_36500[17]}}, p8_bit_slice_36500};
  assign p9_array_37275_comb[12] = {{14{p8_bit_slice_36501[17]}}, p8_bit_slice_36501};
  assign p9_array_37275_comb[13] = {{14{p9_bit_slice_37197_comb[17]}}, p9_bit_slice_37197_comb};
  assign p9_array_37275_comb[14] = {{14{p9_bit_slice_37198_comb[17]}}, p9_bit_slice_37198_comb};
  assign p9_array_37275_comb[15] = {{14{p8_bit_slice_36502[17]}}, p8_bit_slice_36502};
  assign p9_array_37275_comb[16] = {{14{p8_bit_slice_36503[17]}}, p8_bit_slice_36503};
  assign p9_array_37275_comb[17] = {{14{p9_bit_slice_37199_comb[17]}}, p9_bit_slice_37199_comb};
  assign p9_array_37275_comb[18] = {{14{p9_bit_slice_37200_comb[17]}}, p9_bit_slice_37200_comb};
  assign p9_array_37275_comb[19] = {{14{p8_bit_slice_36504[17]}}, p8_bit_slice_36504};
  assign p9_array_37275_comb[20] = {{14{p8_bit_slice_36505[17]}}, p8_bit_slice_36505};
  assign p9_array_37275_comb[21] = {{14{p9_bit_slice_37201_comb[17]}}, p9_bit_slice_37201_comb};
  assign p9_array_37275_comb[22] = {{14{p9_bit_slice_37202_comb[17]}}, p9_bit_slice_37202_comb};
  assign p9_array_37275_comb[23] = {{14{p8_bit_slice_36506[17]}}, p8_bit_slice_36506};
  assign p9_array_37275_comb[24] = {{14{p8_bit_slice_35835[17]}}, p8_bit_slice_35835};
  assign p9_array_37275_comb[25] = {{14{p8_bit_slice_36847[17]}}, p8_bit_slice_36847};
  assign p9_array_37275_comb[26] = {{14{p8_bit_slice_36848[17]}}, p8_bit_slice_36848};
  assign p9_array_37275_comb[27] = {{14{p8_bit_slice_35836[17]}}, p8_bit_slice_35836};
  assign p9_array_37275_comb[28] = {{14{p8_bit_slice_35837[17]}}, p8_bit_slice_35837};
  assign p9_array_37275_comb[29] = {{14{p8_bit_slice_36849[17]}}, p8_bit_slice_36849};
  assign p9_array_37275_comb[30] = {{14{p8_bit_slice_36850[17]}}, p8_bit_slice_36850};
  assign p9_array_37275_comb[31] = {{14{p8_bit_slice_35838[17]}}, p8_bit_slice_35838};
  assign p9_array_37275_comb[32] = {{14{p8_bit_slice_35839[17]}}, p8_bit_slice_35839};
  assign p9_array_37275_comb[33] = {{14{p8_bit_slice_36851[17]}}, p8_bit_slice_36851};
  assign p9_array_37275_comb[34] = {{14{p8_bit_slice_36852[17]}}, p8_bit_slice_36852};
  assign p9_array_37275_comb[35] = {{14{p8_bit_slice_35840[17]}}, p8_bit_slice_35840};
  assign p9_array_37275_comb[36] = {{14{p8_bit_slice_35841[17]}}, p8_bit_slice_35841};
  assign p9_array_37275_comb[37] = {{14{p8_bit_slice_36853[17]}}, p8_bit_slice_36853};
  assign p9_array_37275_comb[38] = {{14{p8_bit_slice_36854[17]}}, p8_bit_slice_36854};
  assign p9_array_37275_comb[39] = {{14{p8_bit_slice_35842[17]}}, p8_bit_slice_35842};
  assign p9_array_37275_comb[40] = {{14{p8_bit_slice_36507[17]}}, p8_bit_slice_36507};
  assign p9_array_37275_comb[41] = {{14{p9_bit_slice_37203_comb[17]}}, p9_bit_slice_37203_comb};
  assign p9_array_37275_comb[42] = {{14{p9_bit_slice_37204_comb[17]}}, p9_bit_slice_37204_comb};
  assign p9_array_37275_comb[43] = {{14{p8_bit_slice_36508[17]}}, p8_bit_slice_36508};
  assign p9_array_37275_comb[44] = {{14{p8_bit_slice_36509[17]}}, p8_bit_slice_36509};
  assign p9_array_37275_comb[45] = {{14{p9_bit_slice_37205_comb[17]}}, p9_bit_slice_37205_comb};
  assign p9_array_37275_comb[46] = {{14{p9_bit_slice_37206_comb[17]}}, p9_bit_slice_37206_comb};
  assign p9_array_37275_comb[47] = {{14{p8_bit_slice_36510[17]}}, p8_bit_slice_36510};
  assign p9_array_37275_comb[48] = {{14{p8_bit_slice_36511[17]}}, p8_bit_slice_36511};
  assign p9_array_37275_comb[49] = {{14{p9_bit_slice_37207_comb[17]}}, p9_bit_slice_37207_comb};
  assign p9_array_37275_comb[50] = {{14{p9_bit_slice_37208_comb[17]}}, p9_bit_slice_37208_comb};
  assign p9_array_37275_comb[51] = {{14{p8_bit_slice_36512[17]}}, p8_bit_slice_36512};
  assign p9_array_37275_comb[52] = {{14{p8_bit_slice_36513[17]}}, p8_bit_slice_36513};
  assign p9_array_37275_comb[53] = {{14{p9_bit_slice_37209_comb[17]}}, p9_bit_slice_37209_comb};
  assign p9_array_37275_comb[54] = {{14{p9_bit_slice_37210_comb[17]}}, p9_bit_slice_37210_comb};
  assign p9_array_37275_comb[55] = {{14{p8_bit_slice_36514[17]}}, p8_bit_slice_36514};
  assign p9_array_37275_comb[56] = {{14{p8_bit_slice_35843[17]}}, p8_bit_slice_35843};
  assign p9_array_37275_comb[57] = {{14{p8_bit_slice_36855[17]}}, p8_bit_slice_36855};
  assign p9_array_37275_comb[58] = {{14{p8_bit_slice_36856[17]}}, p8_bit_slice_36856};
  assign p9_array_37275_comb[59] = {{14{p8_bit_slice_35844[17]}}, p8_bit_slice_35844};
  assign p9_array_37275_comb[60] = {{14{p8_bit_slice_35845[17]}}, p8_bit_slice_35845};
  assign p9_array_37275_comb[61] = {{14{p8_bit_slice_36857[17]}}, p8_bit_slice_36857};
  assign p9_array_37275_comb[62] = {{14{p8_bit_slice_36858[17]}}, p8_bit_slice_36858};
  assign p9_array_37275_comb[63] = {{14{p8_bit_slice_35846[17]}}, p8_bit_slice_35846};

  // Registers for pipe stage 9:
  reg [31:0] p9_array_37275[64];
  always_ff @ (posedge clk) begin
    p9_array_37275 <= p9_array_37275_comb;
  end
  assign out = {p9_array_37275[63], p9_array_37275[62], p9_array_37275[61], p9_array_37275[60], p9_array_37275[59], p9_array_37275[58], p9_array_37275[57], p9_array_37275[56], p9_array_37275[55], p9_array_37275[54], p9_array_37275[53], p9_array_37275[52], p9_array_37275[51], p9_array_37275[50], p9_array_37275[49], p9_array_37275[48], p9_array_37275[47], p9_array_37275[46], p9_array_37275[45], p9_array_37275[44], p9_array_37275[43], p9_array_37275[42], p9_array_37275[41], p9_array_37275[40], p9_array_37275[39], p9_array_37275[38], p9_array_37275[37], p9_array_37275[36], p9_array_37275[35], p9_array_37275[34], p9_array_37275[33], p9_array_37275[32], p9_array_37275[31], p9_array_37275[30], p9_array_37275[29], p9_array_37275[28], p9_array_37275[27], p9_array_37275[26], p9_array_37275[25], p9_array_37275[24], p9_array_37275[23], p9_array_37275[22], p9_array_37275[21], p9_array_37275[20], p9_array_37275[19], p9_array_37275[18], p9_array_37275[17], p9_array_37275[16], p9_array_37275[15], p9_array_37275[14], p9_array_37275[13], p9_array_37275[12], p9_array_37275[11], p9_array_37275[10], p9_array_37275[9], p9_array_37275[8], p9_array_37275[7], p9_array_37275[6], p9_array_37275[5], p9_array_37275[4], p9_array_37275[3], p9_array_37275[2], p9_array_37275[1], p9_array_37275[0]};
endmodule
