module xls_test(
  input wire clk,
  input wire [2047:0] a,
  input wire [2047:0] b,
  input wire [2047:0] result,
  output wire [6143:0] out
);
  // lint_off SIGNED_TYPE
  // lint_off MULTIPLY
  function automatic [31:0] smul32b_32b_x_32b (input reg [31:0] lhs, input reg [31:0] rhs);
    reg signed [31:0] signed_lhs;
    reg signed [31:0] signed_rhs;
    reg signed [31:0] signed_result;
    begin
      signed_lhs = $signed(lhs);
      signed_rhs = $signed(rhs);
      signed_result = signed_lhs * signed_rhs;
      smul32b_32b_x_32b = $unsigned(signed_result);
    end
  endfunction
  // lint_on MULTIPLY
  // lint_on SIGNED_TYPE
  wire [31:0] a_unflattened[8][8];
  assign a_unflattened[0][0] = a[31:0];
  assign a_unflattened[0][1] = a[63:32];
  assign a_unflattened[0][2] = a[95:64];
  assign a_unflattened[0][3] = a[127:96];
  assign a_unflattened[0][4] = a[159:128];
  assign a_unflattened[0][5] = a[191:160];
  assign a_unflattened[0][6] = a[223:192];
  assign a_unflattened[0][7] = a[255:224];
  assign a_unflattened[1][0] = a[287:256];
  assign a_unflattened[1][1] = a[319:288];
  assign a_unflattened[1][2] = a[351:320];
  assign a_unflattened[1][3] = a[383:352];
  assign a_unflattened[1][4] = a[415:384];
  assign a_unflattened[1][5] = a[447:416];
  assign a_unflattened[1][6] = a[479:448];
  assign a_unflattened[1][7] = a[511:480];
  assign a_unflattened[2][0] = a[543:512];
  assign a_unflattened[2][1] = a[575:544];
  assign a_unflattened[2][2] = a[607:576];
  assign a_unflattened[2][3] = a[639:608];
  assign a_unflattened[2][4] = a[671:640];
  assign a_unflattened[2][5] = a[703:672];
  assign a_unflattened[2][6] = a[735:704];
  assign a_unflattened[2][7] = a[767:736];
  assign a_unflattened[3][0] = a[799:768];
  assign a_unflattened[3][1] = a[831:800];
  assign a_unflattened[3][2] = a[863:832];
  assign a_unflattened[3][3] = a[895:864];
  assign a_unflattened[3][4] = a[927:896];
  assign a_unflattened[3][5] = a[959:928];
  assign a_unflattened[3][6] = a[991:960];
  assign a_unflattened[3][7] = a[1023:992];
  assign a_unflattened[4][0] = a[1055:1024];
  assign a_unflattened[4][1] = a[1087:1056];
  assign a_unflattened[4][2] = a[1119:1088];
  assign a_unflattened[4][3] = a[1151:1120];
  assign a_unflattened[4][4] = a[1183:1152];
  assign a_unflattened[4][5] = a[1215:1184];
  assign a_unflattened[4][6] = a[1247:1216];
  assign a_unflattened[4][7] = a[1279:1248];
  assign a_unflattened[5][0] = a[1311:1280];
  assign a_unflattened[5][1] = a[1343:1312];
  assign a_unflattened[5][2] = a[1375:1344];
  assign a_unflattened[5][3] = a[1407:1376];
  assign a_unflattened[5][4] = a[1439:1408];
  assign a_unflattened[5][5] = a[1471:1440];
  assign a_unflattened[5][6] = a[1503:1472];
  assign a_unflattened[5][7] = a[1535:1504];
  assign a_unflattened[6][0] = a[1567:1536];
  assign a_unflattened[6][1] = a[1599:1568];
  assign a_unflattened[6][2] = a[1631:1600];
  assign a_unflattened[6][3] = a[1663:1632];
  assign a_unflattened[6][4] = a[1695:1664];
  assign a_unflattened[6][5] = a[1727:1696];
  assign a_unflattened[6][6] = a[1759:1728];
  assign a_unflattened[6][7] = a[1791:1760];
  assign a_unflattened[7][0] = a[1823:1792];
  assign a_unflattened[7][1] = a[1855:1824];
  assign a_unflattened[7][2] = a[1887:1856];
  assign a_unflattened[7][3] = a[1919:1888];
  assign a_unflattened[7][4] = a[1951:1920];
  assign a_unflattened[7][5] = a[1983:1952];
  assign a_unflattened[7][6] = a[2015:1984];
  assign a_unflattened[7][7] = a[2047:2016];
  wire [31:0] b_unflattened[8][8];
  assign b_unflattened[0][0] = b[31:0];
  assign b_unflattened[0][1] = b[63:32];
  assign b_unflattened[0][2] = b[95:64];
  assign b_unflattened[0][3] = b[127:96];
  assign b_unflattened[0][4] = b[159:128];
  assign b_unflattened[0][5] = b[191:160];
  assign b_unflattened[0][6] = b[223:192];
  assign b_unflattened[0][7] = b[255:224];
  assign b_unflattened[1][0] = b[287:256];
  assign b_unflattened[1][1] = b[319:288];
  assign b_unflattened[1][2] = b[351:320];
  assign b_unflattened[1][3] = b[383:352];
  assign b_unflattened[1][4] = b[415:384];
  assign b_unflattened[1][5] = b[447:416];
  assign b_unflattened[1][6] = b[479:448];
  assign b_unflattened[1][7] = b[511:480];
  assign b_unflattened[2][0] = b[543:512];
  assign b_unflattened[2][1] = b[575:544];
  assign b_unflattened[2][2] = b[607:576];
  assign b_unflattened[2][3] = b[639:608];
  assign b_unflattened[2][4] = b[671:640];
  assign b_unflattened[2][5] = b[703:672];
  assign b_unflattened[2][6] = b[735:704];
  assign b_unflattened[2][7] = b[767:736];
  assign b_unflattened[3][0] = b[799:768];
  assign b_unflattened[3][1] = b[831:800];
  assign b_unflattened[3][2] = b[863:832];
  assign b_unflattened[3][3] = b[895:864];
  assign b_unflattened[3][4] = b[927:896];
  assign b_unflattened[3][5] = b[959:928];
  assign b_unflattened[3][6] = b[991:960];
  assign b_unflattened[3][7] = b[1023:992];
  assign b_unflattened[4][0] = b[1055:1024];
  assign b_unflattened[4][1] = b[1087:1056];
  assign b_unflattened[4][2] = b[1119:1088];
  assign b_unflattened[4][3] = b[1151:1120];
  assign b_unflattened[4][4] = b[1183:1152];
  assign b_unflattened[4][5] = b[1215:1184];
  assign b_unflattened[4][6] = b[1247:1216];
  assign b_unflattened[4][7] = b[1279:1248];
  assign b_unflattened[5][0] = b[1311:1280];
  assign b_unflattened[5][1] = b[1343:1312];
  assign b_unflattened[5][2] = b[1375:1344];
  assign b_unflattened[5][3] = b[1407:1376];
  assign b_unflattened[5][4] = b[1439:1408];
  assign b_unflattened[5][5] = b[1471:1440];
  assign b_unflattened[5][6] = b[1503:1472];
  assign b_unflattened[5][7] = b[1535:1504];
  assign b_unflattened[6][0] = b[1567:1536];
  assign b_unflattened[6][1] = b[1599:1568];
  assign b_unflattened[6][2] = b[1631:1600];
  assign b_unflattened[6][3] = b[1663:1632];
  assign b_unflattened[6][4] = b[1695:1664];
  assign b_unflattened[6][5] = b[1727:1696];
  assign b_unflattened[6][6] = b[1759:1728];
  assign b_unflattened[6][7] = b[1791:1760];
  assign b_unflattened[7][0] = b[1823:1792];
  assign b_unflattened[7][1] = b[1855:1824];
  assign b_unflattened[7][2] = b[1887:1856];
  assign b_unflattened[7][3] = b[1919:1888];
  assign b_unflattened[7][4] = b[1951:1920];
  assign b_unflattened[7][5] = b[1983:1952];
  assign b_unflattened[7][6] = b[2015:1984];
  assign b_unflattened[7][7] = b[2047:2016];
  wire [31:0] result_unflattened[8][8];
  assign result_unflattened[0][0] = result[31:0];
  assign result_unflattened[0][1] = result[63:32];
  assign result_unflattened[0][2] = result[95:64];
  assign result_unflattened[0][3] = result[127:96];
  assign result_unflattened[0][4] = result[159:128];
  assign result_unflattened[0][5] = result[191:160];
  assign result_unflattened[0][6] = result[223:192];
  assign result_unflattened[0][7] = result[255:224];
  assign result_unflattened[1][0] = result[287:256];
  assign result_unflattened[1][1] = result[319:288];
  assign result_unflattened[1][2] = result[351:320];
  assign result_unflattened[1][3] = result[383:352];
  assign result_unflattened[1][4] = result[415:384];
  assign result_unflattened[1][5] = result[447:416];
  assign result_unflattened[1][6] = result[479:448];
  assign result_unflattened[1][7] = result[511:480];
  assign result_unflattened[2][0] = result[543:512];
  assign result_unflattened[2][1] = result[575:544];
  assign result_unflattened[2][2] = result[607:576];
  assign result_unflattened[2][3] = result[639:608];
  assign result_unflattened[2][4] = result[671:640];
  assign result_unflattened[2][5] = result[703:672];
  assign result_unflattened[2][6] = result[735:704];
  assign result_unflattened[2][7] = result[767:736];
  assign result_unflattened[3][0] = result[799:768];
  assign result_unflattened[3][1] = result[831:800];
  assign result_unflattened[3][2] = result[863:832];
  assign result_unflattened[3][3] = result[895:864];
  assign result_unflattened[3][4] = result[927:896];
  assign result_unflattened[3][5] = result[959:928];
  assign result_unflattened[3][6] = result[991:960];
  assign result_unflattened[3][7] = result[1023:992];
  assign result_unflattened[4][0] = result[1055:1024];
  assign result_unflattened[4][1] = result[1087:1056];
  assign result_unflattened[4][2] = result[1119:1088];
  assign result_unflattened[4][3] = result[1151:1120];
  assign result_unflattened[4][4] = result[1183:1152];
  assign result_unflattened[4][5] = result[1215:1184];
  assign result_unflattened[4][6] = result[1247:1216];
  assign result_unflattened[4][7] = result[1279:1248];
  assign result_unflattened[5][0] = result[1311:1280];
  assign result_unflattened[5][1] = result[1343:1312];
  assign result_unflattened[5][2] = result[1375:1344];
  assign result_unflattened[5][3] = result[1407:1376];
  assign result_unflattened[5][4] = result[1439:1408];
  assign result_unflattened[5][5] = result[1471:1440];
  assign result_unflattened[5][6] = result[1503:1472];
  assign result_unflattened[5][7] = result[1535:1504];
  assign result_unflattened[6][0] = result[1567:1536];
  assign result_unflattened[6][1] = result[1599:1568];
  assign result_unflattened[6][2] = result[1631:1600];
  assign result_unflattened[6][3] = result[1663:1632];
  assign result_unflattened[6][4] = result[1695:1664];
  assign result_unflattened[6][5] = result[1727:1696];
  assign result_unflattened[6][6] = result[1759:1728];
  assign result_unflattened[6][7] = result[1791:1760];
  assign result_unflattened[7][0] = result[1823:1792];
  assign result_unflattened[7][1] = result[1855:1824];
  assign result_unflattened[7][2] = result[1887:1856];
  assign result_unflattened[7][3] = result[1919:1888];
  assign result_unflattened[7][4] = result[1951:1920];
  assign result_unflattened[7][5] = result[1983:1952];
  assign result_unflattened[7][6] = result[2015:1984];
  assign result_unflattened[7][7] = result[2047:2016];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_a[8][8];
  reg [31:0] p0_b[8][8];
  always_ff @ (posedge clk) begin
    p0_a <= a_unflattened;
    p0_b <= b_unflattened;
  end

  // ===== Pipe stage 1:
  wire [31:0] p1_array_index_56953_comb;
  wire [31:0] p1_array_index_56954_comb;
  wire [31:0] p1_array_index_56955_comb;
  wire [31:0] p1_array_index_56956_comb;
  wire [31:0] p1_array_index_56961_comb;
  wire [31:0] p1_array_index_56962_comb;
  wire [31:0] p1_array_index_56963_comb;
  wire [31:0] p1_array_index_56964_comb;
  wire [31:0] p1_array_index_56967_comb;
  wire [31:0] p1_array_index_56968_comb;
  wire [31:0] p1_array_index_56971_comb;
  wire [31:0] p1_array_index_56972_comb;
  wire [31:0] p1_array_index_56975_comb;
  wire [31:0] p1_array_index_56976_comb;
  wire [31:0] p1_array_index_56979_comb;
  wire [31:0] p1_array_index_56980_comb;
  wire [31:0] p1_array_index_56983_comb;
  wire [31:0] p1_array_index_56984_comb;
  wire [31:0] p1_array_index_56987_comb;
  wire [31:0] p1_array_index_56988_comb;
  wire [31:0] p1_array_index_56991_comb;
  wire [31:0] p1_array_index_56992_comb;
  wire [31:0] p1_array_index_56995_comb;
  wire [31:0] p1_array_index_56996_comb;
  wire [31:0] p1_array_index_56999_comb;
  wire [31:0] p1_array_index_57000_comb;
  wire [31:0] p1_array_index_57003_comb;
  wire [31:0] p1_array_index_57004_comb;
  wire [31:0] p1_array_index_57007_comb;
  wire [31:0] p1_array_index_57008_comb;
  wire [31:0] p1_array_index_56959_comb;
  wire [31:0] p1_array_index_57011_comb;
  wire [31:0] p1_array_index_56957_comb;
  wire [31:0] p1_array_index_57012_comb;
  wire [31:0] p1_array_index_57015_comb;
  wire [31:0] p1_array_index_57016_comb;
  wire [31:0] p1_array_index_57019_comb;
  wire [31:0] p1_array_index_57020_comb;
  wire [31:0] p1_array_index_57023_comb;
  wire [31:0] p1_array_index_57024_comb;
  wire [31:0] p1_array_index_57027_comb;
  wire [31:0] p1_array_index_57028_comb;
  wire [31:0] p1_array_index_57010_comb;
  wire [31:0] p1_array_index_57009_comb;
  wire [31:0] p1_array_index_57031_comb;
  wire [31:0] p1_array_index_57032_comb;
  wire [31:0] p1_array_index_57035_comb;
  wire [31:0] p1_array_index_57036_comb;
  wire [31:0] p1_array_index_57039_comb;
  wire [31:0] p1_array_index_57040_comb;
  wire [31:0] p1_array_index_57043_comb;
  wire [31:0] p1_array_index_57044_comb;
  wire [31:0] p1_array_index_57047_comb;
  wire [31:0] p1_array_index_57048_comb;
  wire [31:0] p1_array_index_57051_comb;
  wire [31:0] p1_array_index_56960_comb;
  wire [31:0] p1_array_index_57052_comb;
  wire [31:0] p1_array_index_56958_comb;
  wire [31:0] p1_array_index_57050_comb;
  wire [31:0] p1_array_index_57049_comb;
  wire [31:0] p1_array_index_56994_comb;
  wire [31:0] p1_array_index_56993_comb;
  wire [31:0] p1_array_index_57055_comb;
  wire [31:0] p1_array_index_57056_comb;
  wire [31:0] p1_array_index_57059_comb;
  wire [31:0] p1_array_index_57060_comb;
  wire [31:0] p1_array_index_57063_comb;
  wire [31:0] p1_array_index_57064_comb;
  wire [31:0] p1_array_index_57067_comb;
  wire [31:0] p1_array_index_57068_comb;
  wire [31:0] p1_array_index_57071_comb;
  wire [31:0] p1_array_index_57072_comb;
  wire [31:0] p1_array_index_57075_comb;
  wire [31:0] p1_array_index_57076_comb;
  wire [31:0] p1_array_index_57074_comb;
  wire [31:0] p1_array_index_57073_comb;
  wire [31:0] p1_array_index_56951_comb;
  wire [31:0] p1_array_index_56952_comb;
  wire [31:0] p1_array_index_56966_comb;
  wire [31:0] p1_array_index_56970_comb;
  wire [31:0] p1_array_index_56974_comb;
  wire [31:0] p1_array_index_56978_comb;
  wire [31:0] p1_array_index_56982_comb;
  wire [31:0] p1_array_index_56986_comb;
  wire [31:0] p1_array_index_56990_comb;
  wire [31:0] p1_array_index_56998_comb;
  wire [31:0] p1_array_index_57002_comb;
  wire [31:0] p1_array_index_57006_comb;
  wire [31:0] p1_array_index_57014_comb;
  wire [31:0] p1_array_index_57018_comb;
  wire [31:0] p1_array_index_57022_comb;
  wire [31:0] p1_array_index_57026_comb;
  wire [31:0] p1_array_index_57030_comb;
  wire [31:0] p1_array_index_57034_comb;
  wire [31:0] p1_array_index_57038_comb;
  wire [31:0] p1_array_index_57042_comb;
  wire [31:0] p1_array_index_57046_comb;
  wire [31:0] p1_array_index_57054_comb;
  wire [31:0] p1_array_index_57058_comb;
  wire [31:0] p1_array_index_57062_comb;
  wire [31:0] p1_array_index_57066_comb;
  wire [31:0] p1_array_index_57070_comb;
  wire [31:0] p1_array_index_56949_comb;
  wire [31:0] p1_array_index_56950_comb;
  wire [31:0] p1_array_index_56965_comb;
  wire [31:0] p1_array_index_56969_comb;
  wire [31:0] p1_array_index_56973_comb;
  wire [31:0] p1_array_index_56977_comb;
  wire [31:0] p1_array_index_56981_comb;
  wire [31:0] p1_array_index_56985_comb;
  wire [31:0] p1_array_index_56989_comb;
  wire [31:0] p1_array_index_56997_comb;
  wire [31:0] p1_array_index_57001_comb;
  wire [31:0] p1_array_index_57005_comb;
  wire [31:0] p1_array_index_57013_comb;
  wire [31:0] p1_array_index_57017_comb;
  wire [31:0] p1_array_index_57021_comb;
  wire [31:0] p1_array_index_57025_comb;
  wire [31:0] p1_array_index_57029_comb;
  wire [31:0] p1_array_index_57033_comb;
  wire [31:0] p1_array_index_57037_comb;
  wire [31:0] p1_array_index_57041_comb;
  wire [31:0] p1_array_index_57045_comb;
  wire [31:0] p1_array_index_57053_comb;
  wire [31:0] p1_array_index_57057_comb;
  wire [31:0] p1_array_index_57061_comb;
  wire [31:0] p1_array_index_57065_comb;
  wire [31:0] p1_array_index_57069_comb;
  assign p1_array_index_56953_comb = p0_a[3'h0][3'h2];
  assign p1_array_index_56954_comb = p0_b[3'h2][3'h0];
  assign p1_array_index_56955_comb = p0_a[3'h0][3'h3];
  assign p1_array_index_56956_comb = p0_b[3'h3][3'h0];
  assign p1_array_index_56961_comb = p0_a[3'h0][3'h6];
  assign p1_array_index_56962_comb = p0_b[3'h6][3'h0];
  assign p1_array_index_56963_comb = p0_a[3'h0][3'h7];
  assign p1_array_index_56964_comb = p0_b[3'h7][3'h0];
  assign p1_array_index_56967_comb = p0_b[3'h2][3'h1];
  assign p1_array_index_56968_comb = p0_b[3'h3][3'h1];
  assign p1_array_index_56971_comb = p0_b[3'h6][3'h1];
  assign p1_array_index_56972_comb = p0_b[3'h7][3'h1];
  assign p1_array_index_56975_comb = p0_b[3'h2][3'h2];
  assign p1_array_index_56976_comb = p0_b[3'h3][3'h2];
  assign p1_array_index_56979_comb = p0_b[3'h6][3'h2];
  assign p1_array_index_56980_comb = p0_b[3'h7][3'h2];
  assign p1_array_index_56983_comb = p0_b[3'h2][3'h3];
  assign p1_array_index_56984_comb = p0_b[3'h3][3'h3];
  assign p1_array_index_56987_comb = p0_b[3'h6][3'h3];
  assign p1_array_index_56988_comb = p0_b[3'h7][3'h3];
  assign p1_array_index_56991_comb = p0_b[3'h2][3'h4];
  assign p1_array_index_56992_comb = p0_b[3'h3][3'h4];
  assign p1_array_index_56995_comb = p0_b[3'h6][3'h4];
  assign p1_array_index_56996_comb = p0_b[3'h7][3'h4];
  assign p1_array_index_56999_comb = p0_b[3'h2][3'h5];
  assign p1_array_index_57000_comb = p0_b[3'h3][3'h5];
  assign p1_array_index_57003_comb = p0_b[3'h6][3'h5];
  assign p1_array_index_57004_comb = p0_b[3'h7][3'h5];
  assign p1_array_index_57007_comb = p0_b[3'h2][3'h6];
  assign p1_array_index_57008_comb = p0_b[3'h3][3'h6];
  assign p1_array_index_56959_comb = p0_a[3'h0][3'h4];
  assign p1_array_index_57011_comb = p0_b[3'h4][3'h6];
  assign p1_array_index_56957_comb = p0_a[3'h0][3'h5];
  assign p1_array_index_57012_comb = p0_b[3'h5][3'h6];
  assign p1_array_index_57015_comb = p0_b[3'h2][3'h7];
  assign p1_array_index_57016_comb = p0_b[3'h3][3'h7];
  assign p1_array_index_57019_comb = p0_b[3'h6][3'h7];
  assign p1_array_index_57020_comb = p0_b[3'h7][3'h7];
  assign p1_array_index_57023_comb = p0_a[3'h1][3'h2];
  assign p1_array_index_57024_comb = p0_a[3'h1][3'h3];
  assign p1_array_index_57027_comb = p0_a[3'h1][3'h6];
  assign p1_array_index_57028_comb = p0_a[3'h1][3'h7];
  assign p1_array_index_57010_comb = p0_b[3'h6][3'h6];
  assign p1_array_index_57009_comb = p0_b[3'h7][3'h6];
  assign p1_array_index_57031_comb = p0_a[3'h2][3'h2];
  assign p1_array_index_57032_comb = p0_a[3'h2][3'h3];
  assign p1_array_index_57035_comb = p0_a[3'h2][3'h6];
  assign p1_array_index_57036_comb = p0_a[3'h2][3'h7];
  assign p1_array_index_57039_comb = p0_a[3'h3][3'h2];
  assign p1_array_index_57040_comb = p0_a[3'h3][3'h3];
  assign p1_array_index_57043_comb = p0_a[3'h3][3'h6];
  assign p1_array_index_57044_comb = p0_a[3'h3][3'h7];
  assign p1_array_index_57047_comb = p0_a[3'h4][3'h2];
  assign p1_array_index_57048_comb = p0_a[3'h4][3'h3];
  assign p1_array_index_57051_comb = p0_a[3'h4][3'h4];
  assign p1_array_index_56960_comb = p0_b[3'h4][3'h0];
  assign p1_array_index_57052_comb = p0_a[3'h4][3'h5];
  assign p1_array_index_56958_comb = p0_b[3'h5][3'h0];
  assign p1_array_index_57050_comb = p0_a[3'h4][3'h6];
  assign p1_array_index_57049_comb = p0_a[3'h4][3'h7];
  assign p1_array_index_56994_comb = p0_b[3'h4][3'h4];
  assign p1_array_index_56993_comb = p0_b[3'h5][3'h4];
  assign p1_array_index_57055_comb = p0_a[3'h5][3'h2];
  assign p1_array_index_57056_comb = p0_a[3'h5][3'h3];
  assign p1_array_index_57059_comb = p0_a[3'h5][3'h6];
  assign p1_array_index_57060_comb = p0_a[3'h5][3'h7];
  assign p1_array_index_57063_comb = p0_a[3'h6][3'h2];
  assign p1_array_index_57064_comb = p0_a[3'h6][3'h3];
  assign p1_array_index_57067_comb = p0_a[3'h6][3'h6];
  assign p1_array_index_57068_comb = p0_a[3'h6][3'h7];
  assign p1_array_index_57071_comb = p0_a[3'h7][3'h2];
  assign p1_array_index_57072_comb = p0_a[3'h7][3'h3];
  assign p1_array_index_57075_comb = p0_a[3'h7][3'h4];
  assign p1_array_index_57076_comb = p0_a[3'h7][3'h5];
  assign p1_array_index_57074_comb = p0_a[3'h7][3'h6];
  assign p1_array_index_57073_comb = p0_a[3'h7][3'h7];
  assign p1_array_index_56951_comb = p0_a[3'h0][3'h0];
  assign p1_array_index_56952_comb = p0_b[3'h0][3'h0];
  assign p1_array_index_56966_comb = p0_b[3'h0][3'h1];
  assign p1_array_index_56970_comb = p0_b[3'h4][3'h1];
  assign p1_array_index_56974_comb = p0_b[3'h0][3'h2];
  assign p1_array_index_56978_comb = p0_b[3'h4][3'h2];
  assign p1_array_index_56982_comb = p0_b[3'h0][3'h3];
  assign p1_array_index_56986_comb = p0_b[3'h4][3'h3];
  assign p1_array_index_56990_comb = p0_b[3'h0][3'h4];
  assign p1_array_index_56998_comb = p0_b[3'h0][3'h5];
  assign p1_array_index_57002_comb = p0_b[3'h4][3'h5];
  assign p1_array_index_57006_comb = p0_b[3'h0][3'h6];
  assign p1_array_index_57014_comb = p0_b[3'h0][3'h7];
  assign p1_array_index_57018_comb = p0_b[3'h4][3'h7];
  assign p1_array_index_57022_comb = p0_a[3'h1][3'h0];
  assign p1_array_index_57026_comb = p0_a[3'h1][3'h4];
  assign p1_array_index_57030_comb = p0_a[3'h2][3'h0];
  assign p1_array_index_57034_comb = p0_a[3'h2][3'h4];
  assign p1_array_index_57038_comb = p0_a[3'h3][3'h0];
  assign p1_array_index_57042_comb = p0_a[3'h3][3'h4];
  assign p1_array_index_57046_comb = p0_a[3'h4][3'h0];
  assign p1_array_index_57054_comb = p0_a[3'h5][3'h0];
  assign p1_array_index_57058_comb = p0_a[3'h5][3'h4];
  assign p1_array_index_57062_comb = p0_a[3'h6][3'h0];
  assign p1_array_index_57066_comb = p0_a[3'h6][3'h4];
  assign p1_array_index_57070_comb = p0_a[3'h7][3'h0];
  assign p1_array_index_56949_comb = p0_a[3'h0][3'h1];
  assign p1_array_index_56950_comb = p0_b[3'h1][3'h0];
  assign p1_array_index_56965_comb = p0_b[3'h1][3'h1];
  assign p1_array_index_56969_comb = p0_b[3'h5][3'h1];
  assign p1_array_index_56973_comb = p0_b[3'h1][3'h2];
  assign p1_array_index_56977_comb = p0_b[3'h5][3'h2];
  assign p1_array_index_56981_comb = p0_b[3'h1][3'h3];
  assign p1_array_index_56985_comb = p0_b[3'h5][3'h3];
  assign p1_array_index_56989_comb = p0_b[3'h1][3'h4];
  assign p1_array_index_56997_comb = p0_b[3'h1][3'h5];
  assign p1_array_index_57001_comb = p0_b[3'h5][3'h5];
  assign p1_array_index_57005_comb = p0_b[3'h1][3'h6];
  assign p1_array_index_57013_comb = p0_b[3'h1][3'h7];
  assign p1_array_index_57017_comb = p0_b[3'h5][3'h7];
  assign p1_array_index_57021_comb = p0_a[3'h1][3'h1];
  assign p1_array_index_57025_comb = p0_a[3'h1][3'h5];
  assign p1_array_index_57029_comb = p0_a[3'h2][3'h1];
  assign p1_array_index_57033_comb = p0_a[3'h2][3'h5];
  assign p1_array_index_57037_comb = p0_a[3'h3][3'h1];
  assign p1_array_index_57041_comb = p0_a[3'h3][3'h5];
  assign p1_array_index_57045_comb = p0_a[3'h4][3'h1];
  assign p1_array_index_57053_comb = p0_a[3'h5][3'h1];
  assign p1_array_index_57057_comb = p0_a[3'h5][3'h5];
  assign p1_array_index_57061_comb = p0_a[3'h6][3'h1];
  assign p1_array_index_57065_comb = p0_a[3'h6][3'h5];
  assign p1_array_index_57069_comb = p0_a[3'h7][3'h1];

  // Registers for pipe stage 1:
  reg [31:0] p1_a[8][8];
  reg [31:0] p1_b[8][8];
  reg [31:0] p1_array_index_56953;
  reg [31:0] p1_array_index_56954;
  reg [31:0] p1_array_index_56955;
  reg [31:0] p1_array_index_56956;
  reg [31:0] p1_array_index_56961;
  reg [31:0] p1_array_index_56962;
  reg [31:0] p1_array_index_56963;
  reg [31:0] p1_array_index_56964;
  reg [31:0] p1_array_index_56967;
  reg [31:0] p1_array_index_56968;
  reg [31:0] p1_array_index_56971;
  reg [31:0] p1_array_index_56972;
  reg [31:0] p1_array_index_56975;
  reg [31:0] p1_array_index_56976;
  reg [31:0] p1_array_index_56979;
  reg [31:0] p1_array_index_56980;
  reg [31:0] p1_array_index_56983;
  reg [31:0] p1_array_index_56984;
  reg [31:0] p1_array_index_56987;
  reg [31:0] p1_array_index_56988;
  reg [31:0] p1_array_index_56991;
  reg [31:0] p1_array_index_56992;
  reg [31:0] p1_array_index_56995;
  reg [31:0] p1_array_index_56996;
  reg [31:0] p1_array_index_56999;
  reg [31:0] p1_array_index_57000;
  reg [31:0] p1_array_index_57003;
  reg [31:0] p1_array_index_57004;
  reg [31:0] p1_array_index_57007;
  reg [31:0] p1_array_index_57008;
  reg [31:0] p1_array_index_56959;
  reg [31:0] p1_array_index_57011;
  reg [31:0] p1_array_index_56957;
  reg [31:0] p1_array_index_57012;
  reg [31:0] p1_array_index_57015;
  reg [31:0] p1_array_index_57016;
  reg [31:0] p1_array_index_57019;
  reg [31:0] p1_array_index_57020;
  reg [31:0] p1_array_index_57023;
  reg [31:0] p1_array_index_57024;
  reg [31:0] p1_array_index_57027;
  reg [31:0] p1_array_index_57028;
  reg [31:0] p1_array_index_57010;
  reg [31:0] p1_array_index_57009;
  reg [31:0] p1_array_index_57031;
  reg [31:0] p1_array_index_57032;
  reg [31:0] p1_array_index_57035;
  reg [31:0] p1_array_index_57036;
  reg [31:0] p1_array_index_57039;
  reg [31:0] p1_array_index_57040;
  reg [31:0] p1_array_index_57043;
  reg [31:0] p1_array_index_57044;
  reg [31:0] p1_array_index_57047;
  reg [31:0] p1_array_index_57048;
  reg [31:0] p1_array_index_57051;
  reg [31:0] p1_array_index_56960;
  reg [31:0] p1_array_index_57052;
  reg [31:0] p1_array_index_56958;
  reg [31:0] p1_array_index_57050;
  reg [31:0] p1_array_index_57049;
  reg [31:0] p1_array_index_56994;
  reg [31:0] p1_array_index_56993;
  reg [31:0] p1_array_index_57055;
  reg [31:0] p1_array_index_57056;
  reg [31:0] p1_array_index_57059;
  reg [31:0] p1_array_index_57060;
  reg [31:0] p1_array_index_57063;
  reg [31:0] p1_array_index_57064;
  reg [31:0] p1_array_index_57067;
  reg [31:0] p1_array_index_57068;
  reg [31:0] p1_array_index_57071;
  reg [31:0] p1_array_index_57072;
  reg [31:0] p1_array_index_57075;
  reg [31:0] p1_array_index_57076;
  reg [31:0] p1_array_index_57074;
  reg [31:0] p1_array_index_57073;
  reg [31:0] p1_array_index_56951;
  reg [31:0] p1_array_index_56952;
  reg [31:0] p1_array_index_56966;
  reg [31:0] p1_array_index_56970;
  reg [31:0] p1_array_index_56974;
  reg [31:0] p1_array_index_56978;
  reg [31:0] p1_array_index_56982;
  reg [31:0] p1_array_index_56986;
  reg [31:0] p1_array_index_56990;
  reg [31:0] p1_array_index_56998;
  reg [31:0] p1_array_index_57002;
  reg [31:0] p1_array_index_57006;
  reg [31:0] p1_array_index_57014;
  reg [31:0] p1_array_index_57018;
  reg [31:0] p1_array_index_57022;
  reg [31:0] p1_array_index_57026;
  reg [31:0] p1_array_index_57030;
  reg [31:0] p1_array_index_57034;
  reg [31:0] p1_array_index_57038;
  reg [31:0] p1_array_index_57042;
  reg [31:0] p1_array_index_57046;
  reg [31:0] p1_array_index_57054;
  reg [31:0] p1_array_index_57058;
  reg [31:0] p1_array_index_57062;
  reg [31:0] p1_array_index_57066;
  reg [31:0] p1_array_index_57070;
  reg [31:0] p1_array_index_56949;
  reg [31:0] p1_array_index_56950;
  reg [31:0] p1_array_index_56965;
  reg [31:0] p1_array_index_56969;
  reg [31:0] p1_array_index_56973;
  reg [31:0] p1_array_index_56977;
  reg [31:0] p1_array_index_56981;
  reg [31:0] p1_array_index_56985;
  reg [31:0] p1_array_index_56989;
  reg [31:0] p1_array_index_56997;
  reg [31:0] p1_array_index_57001;
  reg [31:0] p1_array_index_57005;
  reg [31:0] p1_array_index_57013;
  reg [31:0] p1_array_index_57017;
  reg [31:0] p1_array_index_57021;
  reg [31:0] p1_array_index_57025;
  reg [31:0] p1_array_index_57029;
  reg [31:0] p1_array_index_57033;
  reg [31:0] p1_array_index_57037;
  reg [31:0] p1_array_index_57041;
  reg [31:0] p1_array_index_57045;
  reg [31:0] p1_array_index_57053;
  reg [31:0] p1_array_index_57057;
  reg [31:0] p1_array_index_57061;
  reg [31:0] p1_array_index_57065;
  reg [31:0] p1_array_index_57069;
  always_ff @ (posedge clk) begin
    p1_a <= p0_a;
    p1_b <= p0_b;
    p1_array_index_56953 <= p1_array_index_56953_comb;
    p1_array_index_56954 <= p1_array_index_56954_comb;
    p1_array_index_56955 <= p1_array_index_56955_comb;
    p1_array_index_56956 <= p1_array_index_56956_comb;
    p1_array_index_56961 <= p1_array_index_56961_comb;
    p1_array_index_56962 <= p1_array_index_56962_comb;
    p1_array_index_56963 <= p1_array_index_56963_comb;
    p1_array_index_56964 <= p1_array_index_56964_comb;
    p1_array_index_56967 <= p1_array_index_56967_comb;
    p1_array_index_56968 <= p1_array_index_56968_comb;
    p1_array_index_56971 <= p1_array_index_56971_comb;
    p1_array_index_56972 <= p1_array_index_56972_comb;
    p1_array_index_56975 <= p1_array_index_56975_comb;
    p1_array_index_56976 <= p1_array_index_56976_comb;
    p1_array_index_56979 <= p1_array_index_56979_comb;
    p1_array_index_56980 <= p1_array_index_56980_comb;
    p1_array_index_56983 <= p1_array_index_56983_comb;
    p1_array_index_56984 <= p1_array_index_56984_comb;
    p1_array_index_56987 <= p1_array_index_56987_comb;
    p1_array_index_56988 <= p1_array_index_56988_comb;
    p1_array_index_56991 <= p1_array_index_56991_comb;
    p1_array_index_56992 <= p1_array_index_56992_comb;
    p1_array_index_56995 <= p1_array_index_56995_comb;
    p1_array_index_56996 <= p1_array_index_56996_comb;
    p1_array_index_56999 <= p1_array_index_56999_comb;
    p1_array_index_57000 <= p1_array_index_57000_comb;
    p1_array_index_57003 <= p1_array_index_57003_comb;
    p1_array_index_57004 <= p1_array_index_57004_comb;
    p1_array_index_57007 <= p1_array_index_57007_comb;
    p1_array_index_57008 <= p1_array_index_57008_comb;
    p1_array_index_56959 <= p1_array_index_56959_comb;
    p1_array_index_57011 <= p1_array_index_57011_comb;
    p1_array_index_56957 <= p1_array_index_56957_comb;
    p1_array_index_57012 <= p1_array_index_57012_comb;
    p1_array_index_57015 <= p1_array_index_57015_comb;
    p1_array_index_57016 <= p1_array_index_57016_comb;
    p1_array_index_57019 <= p1_array_index_57019_comb;
    p1_array_index_57020 <= p1_array_index_57020_comb;
    p1_array_index_57023 <= p1_array_index_57023_comb;
    p1_array_index_57024 <= p1_array_index_57024_comb;
    p1_array_index_57027 <= p1_array_index_57027_comb;
    p1_array_index_57028 <= p1_array_index_57028_comb;
    p1_array_index_57010 <= p1_array_index_57010_comb;
    p1_array_index_57009 <= p1_array_index_57009_comb;
    p1_array_index_57031 <= p1_array_index_57031_comb;
    p1_array_index_57032 <= p1_array_index_57032_comb;
    p1_array_index_57035 <= p1_array_index_57035_comb;
    p1_array_index_57036 <= p1_array_index_57036_comb;
    p1_array_index_57039 <= p1_array_index_57039_comb;
    p1_array_index_57040 <= p1_array_index_57040_comb;
    p1_array_index_57043 <= p1_array_index_57043_comb;
    p1_array_index_57044 <= p1_array_index_57044_comb;
    p1_array_index_57047 <= p1_array_index_57047_comb;
    p1_array_index_57048 <= p1_array_index_57048_comb;
    p1_array_index_57051 <= p1_array_index_57051_comb;
    p1_array_index_56960 <= p1_array_index_56960_comb;
    p1_array_index_57052 <= p1_array_index_57052_comb;
    p1_array_index_56958 <= p1_array_index_56958_comb;
    p1_array_index_57050 <= p1_array_index_57050_comb;
    p1_array_index_57049 <= p1_array_index_57049_comb;
    p1_array_index_56994 <= p1_array_index_56994_comb;
    p1_array_index_56993 <= p1_array_index_56993_comb;
    p1_array_index_57055 <= p1_array_index_57055_comb;
    p1_array_index_57056 <= p1_array_index_57056_comb;
    p1_array_index_57059 <= p1_array_index_57059_comb;
    p1_array_index_57060 <= p1_array_index_57060_comb;
    p1_array_index_57063 <= p1_array_index_57063_comb;
    p1_array_index_57064 <= p1_array_index_57064_comb;
    p1_array_index_57067 <= p1_array_index_57067_comb;
    p1_array_index_57068 <= p1_array_index_57068_comb;
    p1_array_index_57071 <= p1_array_index_57071_comb;
    p1_array_index_57072 <= p1_array_index_57072_comb;
    p1_array_index_57075 <= p1_array_index_57075_comb;
    p1_array_index_57076 <= p1_array_index_57076_comb;
    p1_array_index_57074 <= p1_array_index_57074_comb;
    p1_array_index_57073 <= p1_array_index_57073_comb;
    p1_array_index_56951 <= p1_array_index_56951_comb;
    p1_array_index_56952 <= p1_array_index_56952_comb;
    p1_array_index_56966 <= p1_array_index_56966_comb;
    p1_array_index_56970 <= p1_array_index_56970_comb;
    p1_array_index_56974 <= p1_array_index_56974_comb;
    p1_array_index_56978 <= p1_array_index_56978_comb;
    p1_array_index_56982 <= p1_array_index_56982_comb;
    p1_array_index_56986 <= p1_array_index_56986_comb;
    p1_array_index_56990 <= p1_array_index_56990_comb;
    p1_array_index_56998 <= p1_array_index_56998_comb;
    p1_array_index_57002 <= p1_array_index_57002_comb;
    p1_array_index_57006 <= p1_array_index_57006_comb;
    p1_array_index_57014 <= p1_array_index_57014_comb;
    p1_array_index_57018 <= p1_array_index_57018_comb;
    p1_array_index_57022 <= p1_array_index_57022_comb;
    p1_array_index_57026 <= p1_array_index_57026_comb;
    p1_array_index_57030 <= p1_array_index_57030_comb;
    p1_array_index_57034 <= p1_array_index_57034_comb;
    p1_array_index_57038 <= p1_array_index_57038_comb;
    p1_array_index_57042 <= p1_array_index_57042_comb;
    p1_array_index_57046 <= p1_array_index_57046_comb;
    p1_array_index_57054 <= p1_array_index_57054_comb;
    p1_array_index_57058 <= p1_array_index_57058_comb;
    p1_array_index_57062 <= p1_array_index_57062_comb;
    p1_array_index_57066 <= p1_array_index_57066_comb;
    p1_array_index_57070 <= p1_array_index_57070_comb;
    p1_array_index_56949 <= p1_array_index_56949_comb;
    p1_array_index_56950 <= p1_array_index_56950_comb;
    p1_array_index_56965 <= p1_array_index_56965_comb;
    p1_array_index_56969 <= p1_array_index_56969_comb;
    p1_array_index_56973 <= p1_array_index_56973_comb;
    p1_array_index_56977 <= p1_array_index_56977_comb;
    p1_array_index_56981 <= p1_array_index_56981_comb;
    p1_array_index_56985 <= p1_array_index_56985_comb;
    p1_array_index_56989 <= p1_array_index_56989_comb;
    p1_array_index_56997 <= p1_array_index_56997_comb;
    p1_array_index_57001 <= p1_array_index_57001_comb;
    p1_array_index_57005 <= p1_array_index_57005_comb;
    p1_array_index_57013 <= p1_array_index_57013_comb;
    p1_array_index_57017 <= p1_array_index_57017_comb;
    p1_array_index_57021 <= p1_array_index_57021_comb;
    p1_array_index_57025 <= p1_array_index_57025_comb;
    p1_array_index_57029 <= p1_array_index_57029_comb;
    p1_array_index_57033 <= p1_array_index_57033_comb;
    p1_array_index_57037 <= p1_array_index_57037_comb;
    p1_array_index_57041 <= p1_array_index_57041_comb;
    p1_array_index_57045 <= p1_array_index_57045_comb;
    p1_array_index_57053 <= p1_array_index_57053_comb;
    p1_array_index_57057 <= p1_array_index_57057_comb;
    p1_array_index_57061 <= p1_array_index_57061_comb;
    p1_array_index_57065 <= p1_array_index_57065_comb;
    p1_array_index_57069 <= p1_array_index_57069_comb;
  end

  // ===== Pipe stage 2:
  wire [31:0] p2_smul_57841_comb;
  wire [31:0] p2_smul_57842_comb;
  wire [31:0] p2_smul_57843_comb;
  wire [31:0] p2_smul_57844_comb;
  wire [31:0] p2_smul_57845_comb;
  wire [31:0] p2_smul_57846_comb;
  wire [31:0] p2_smul_57847_comb;
  wire [31:0] p2_smul_57848_comb;
  wire [31:0] p2_smul_57833_comb;
  wire [31:0] p2_smul_57834_comb;
  wire [31:0] p2_smul_57835_comb;
  wire [31:0] p2_smul_57836_comb;
  wire [31:0] p2_smul_57837_comb;
  wire [31:0] p2_smul_57838_comb;
  wire [31:0] p2_smul_57839_comb;
  wire [31:0] p2_smul_57840_comb;
  wire [31:0] p2_smul_57825_comb;
  wire [31:0] p2_smul_57826_comb;
  wire [31:0] p2_smul_57827_comb;
  wire [31:0] p2_smul_57828_comb;
  wire [31:0] p2_smul_57829_comb;
  wire [31:0] p2_smul_57830_comb;
  wire [31:0] p2_smul_57831_comb;
  wire [31:0] p2_smul_57832_comb;
  wire [31:0] p2_smul_57817_comb;
  wire [31:0] p2_smul_57818_comb;
  wire [31:0] p2_smul_57819_comb;
  wire [31:0] p2_smul_57820_comb;
  wire [31:0] p2_smul_57821_comb;
  wire [31:0] p2_smul_57822_comb;
  wire [31:0] p2_smul_57823_comb;
  wire [31:0] p2_smul_57824_comb;
  wire [31:0] p2_smul_57809_comb;
  wire [31:0] p2_smul_57810_comb;
  wire [31:0] p2_smul_57811_comb;
  wire [31:0] p2_smul_57812_comb;
  wire [31:0] p2_smul_57813_comb;
  wire [31:0] p2_smul_57814_comb;
  wire [31:0] p2_smul_57815_comb;
  wire [31:0] p2_smul_57816_comb;
  wire [31:0] p2_smul_57801_comb;
  wire [31:0] p2_smul_57802_comb;
  wire [31:0] p2_smul_57803_comb;
  wire [31:0] p2_smul_57804_comb;
  wire [31:0] p2_smul_57805_comb;
  wire [31:0] p2_smul_57806_comb;
  wire [31:0] p2_smul_57807_comb;
  wire [31:0] p2_smul_57808_comb;
  wire [31:0] p2_smul_57793_comb;
  wire [31:0] p2_smul_57794_comb;
  wire [31:0] p2_smul_57795_comb;
  wire [31:0] p2_smul_57796_comb;
  wire [31:0] p2_smul_57797_comb;
  wire [31:0] p2_smul_57798_comb;
  wire [31:0] p2_smul_57799_comb;
  wire [31:0] p2_smul_57800_comb;
  wire [31:0] p2_smul_57785_comb;
  wire [31:0] p2_smul_57786_comb;
  wire [31:0] p2_smul_57787_comb;
  wire [31:0] p2_smul_57788_comb;
  wire [31:0] p2_smul_57789_comb;
  wire [31:0] p2_smul_57790_comb;
  wire [31:0] p2_smul_57791_comb;
  wire [31:0] p2_smul_57792_comb;
  wire [31:0] p2_smul_57777_comb;
  wire [31:0] p2_smul_57778_comb;
  wire [31:0] p2_smul_57779_comb;
  wire [31:0] p2_smul_57780_comb;
  wire [31:0] p2_smul_57781_comb;
  wire [31:0] p2_smul_57782_comb;
  wire [31:0] p2_smul_57783_comb;
  wire [31:0] p2_smul_57784_comb;
  wire [31:0] p2_smul_57769_comb;
  wire [31:0] p2_smul_57770_comb;
  wire [31:0] p2_smul_57771_comb;
  wire [31:0] p2_smul_57772_comb;
  wire [31:0] p2_smul_57773_comb;
  wire [31:0] p2_smul_57774_comb;
  wire [31:0] p2_smul_57775_comb;
  wire [31:0] p2_smul_57776_comb;
  wire [31:0] p2_smul_57761_comb;
  wire [31:0] p2_smul_57762_comb;
  wire [31:0] p2_smul_57763_comb;
  wire [31:0] p2_smul_57764_comb;
  wire [31:0] p2_smul_57765_comb;
  wire [31:0] p2_smul_57766_comb;
  wire [31:0] p2_smul_57767_comb;
  wire [31:0] p2_smul_57768_comb;
  wire [31:0] p2_smul_57753_comb;
  wire [31:0] p2_smul_57754_comb;
  wire [31:0] p2_smul_57755_comb;
  wire [31:0] p2_smul_57756_comb;
  wire [31:0] p2_smul_57757_comb;
  wire [31:0] p2_smul_57758_comb;
  wire [31:0] p2_smul_57759_comb;
  wire [31:0] p2_smul_57760_comb;
  wire [31:0] p2_smul_57745_comb;
  wire [31:0] p2_smul_57746_comb;
  wire [31:0] p2_smul_57747_comb;
  wire [31:0] p2_smul_57748_comb;
  wire [31:0] p2_smul_57749_comb;
  wire [31:0] p2_smul_57750_comb;
  wire [31:0] p2_smul_57751_comb;
  wire [31:0] p2_smul_57752_comb;
  wire [31:0] p2_smul_57737_comb;
  wire [31:0] p2_smul_57738_comb;
  wire [31:0] p2_smul_57739_comb;
  wire [31:0] p2_smul_57740_comb;
  wire [31:0] p2_smul_57741_comb;
  wire [31:0] p2_smul_57742_comb;
  wire [31:0] p2_smul_57743_comb;
  wire [31:0] p2_smul_57744_comb;
  wire [31:0] p2_smul_57729_comb;
  wire [31:0] p2_smul_57730_comb;
  wire [31:0] p2_smul_57731_comb;
  wire [31:0] p2_smul_57732_comb;
  wire [31:0] p2_smul_57733_comb;
  wire [31:0] p2_smul_57734_comb;
  wire [31:0] p2_smul_57735_comb;
  wire [31:0] p2_smul_57736_comb;
  wire [31:0] p2_smul_57721_comb;
  wire [31:0] p2_smul_57722_comb;
  wire [31:0] p2_smul_57723_comb;
  wire [31:0] p2_smul_57724_comb;
  wire [31:0] p2_smul_57725_comb;
  wire [31:0] p2_smul_57726_comb;
  wire [31:0] p2_smul_57727_comb;
  wire [31:0] p2_smul_57728_comb;
  wire [31:0] p2_smul_57713_comb;
  wire [31:0] p2_smul_57714_comb;
  wire [31:0] p2_smul_57715_comb;
  wire [31:0] p2_smul_57716_comb;
  wire [31:0] p2_smul_57717_comb;
  wire [31:0] p2_smul_57718_comb;
  wire [31:0] p2_smul_57719_comb;
  wire [31:0] p2_smul_57720_comb;
  wire [31:0] p2_smul_57705_comb;
  wire [31:0] p2_smul_57706_comb;
  wire [31:0] p2_smul_57707_comb;
  wire [31:0] p2_smul_57708_comb;
  wire [31:0] p2_smul_57709_comb;
  wire [31:0] p2_smul_57710_comb;
  wire [31:0] p2_smul_57711_comb;
  wire [31:0] p2_smul_57712_comb;
  wire [31:0] p2_smul_57697_comb;
  wire [31:0] p2_smul_57698_comb;
  wire [31:0] p2_smul_57699_comb;
  wire [31:0] p2_smul_57700_comb;
  wire [31:0] p2_smul_57701_comb;
  wire [31:0] p2_smul_57702_comb;
  wire [31:0] p2_smul_57703_comb;
  wire [31:0] p2_smul_57704_comb;
  wire [31:0] p2_smul_57689_comb;
  wire [31:0] p2_smul_57690_comb;
  wire [31:0] p2_smul_57691_comb;
  wire [31:0] p2_smul_57692_comb;
  wire [31:0] p2_smul_57693_comb;
  wire [31:0] p2_smul_57694_comb;
  wire [31:0] p2_smul_57695_comb;
  wire [31:0] p2_smul_57696_comb;
  wire [31:0] p2_smul_57681_comb;
  wire [31:0] p2_smul_57682_comb;
  wire [31:0] p2_smul_57683_comb;
  wire [31:0] p2_smul_57684_comb;
  wire [31:0] p2_smul_57685_comb;
  wire [31:0] p2_smul_57686_comb;
  wire [31:0] p2_smul_57687_comb;
  wire [31:0] p2_smul_57688_comb;
  wire [31:0] p2_smul_57673_comb;
  wire [31:0] p2_smul_57674_comb;
  wire [31:0] p2_smul_57675_comb;
  wire [31:0] p2_smul_57676_comb;
  wire [31:0] p2_smul_57677_comb;
  wire [31:0] p2_smul_57678_comb;
  wire [31:0] p2_smul_57679_comb;
  wire [31:0] p2_smul_57680_comb;
  wire [31:0] p2_smul_57665_comb;
  wire [31:0] p2_smul_57666_comb;
  wire [31:0] p2_smul_57667_comb;
  wire [31:0] p2_smul_57668_comb;
  wire [31:0] p2_smul_57669_comb;
  wire [31:0] p2_smul_57670_comb;
  wire [31:0] p2_smul_57671_comb;
  wire [31:0] p2_smul_57672_comb;
  wire [31:0] p2_smul_57657_comb;
  wire [31:0] p2_smul_57658_comb;
  wire [31:0] p2_smul_57659_comb;
  wire [31:0] p2_smul_57660_comb;
  wire [31:0] p2_smul_57661_comb;
  wire [31:0] p2_smul_57662_comb;
  wire [31:0] p2_smul_57663_comb;
  wire [31:0] p2_smul_57664_comb;
  wire [31:0] p2_smul_57649_comb;
  wire [31:0] p2_smul_57650_comb;
  wire [31:0] p2_smul_57651_comb;
  wire [31:0] p2_smul_57652_comb;
  wire [31:0] p2_smul_57653_comb;
  wire [31:0] p2_smul_57654_comb;
  wire [31:0] p2_smul_57655_comb;
  wire [31:0] p2_smul_57656_comb;
  wire [31:0] p2_smul_57641_comb;
  wire [31:0] p2_smul_57642_comb;
  wire [31:0] p2_smul_57643_comb;
  wire [31:0] p2_smul_57644_comb;
  wire [31:0] p2_smul_57645_comb;
  wire [31:0] p2_smul_57646_comb;
  wire [31:0] p2_smul_57647_comb;
  wire [31:0] p2_smul_57648_comb;
  wire [31:0] p2_smul_57633_comb;
  wire [31:0] p2_smul_57634_comb;
  wire [31:0] p2_smul_57635_comb;
  wire [31:0] p2_smul_57636_comb;
  wire [31:0] p2_smul_57637_comb;
  wire [31:0] p2_smul_57638_comb;
  wire [31:0] p2_smul_57639_comb;
  wire [31:0] p2_smul_57640_comb;
  wire [31:0] p2_smul_57625_comb;
  wire [31:0] p2_smul_57626_comb;
  wire [31:0] p2_smul_57627_comb;
  wire [31:0] p2_smul_57628_comb;
  wire [31:0] p2_smul_57629_comb;
  wire [31:0] p2_smul_57630_comb;
  wire [31:0] p2_smul_57631_comb;
  wire [31:0] p2_smul_57632_comb;
  wire [31:0] p2_smul_57617_comb;
  wire [31:0] p2_smul_57618_comb;
  wire [31:0] p2_smul_57619_comb;
  wire [31:0] p2_smul_57620_comb;
  wire [31:0] p2_smul_57621_comb;
  wire [31:0] p2_smul_57622_comb;
  wire [31:0] p2_smul_57623_comb;
  wire [31:0] p2_smul_57624_comb;
  wire [31:0] p2_smul_57609_comb;
  wire [31:0] p2_smul_57610_comb;
  wire [31:0] p2_smul_57611_comb;
  wire [31:0] p2_smul_57612_comb;
  wire [31:0] p2_smul_57613_comb;
  wire [31:0] p2_smul_57614_comb;
  wire [31:0] p2_smul_57615_comb;
  wire [31:0] p2_smul_57616_comb;
  wire [31:0] p2_smul_57601_comb;
  wire [31:0] p2_smul_57602_comb;
  wire [31:0] p2_smul_57603_comb;
  wire [31:0] p2_smul_57604_comb;
  wire [31:0] p2_smul_57605_comb;
  wire [31:0] p2_smul_57606_comb;
  wire [31:0] p2_smul_57607_comb;
  wire [31:0] p2_smul_57608_comb;
  wire [31:0] p2_smul_57593_comb;
  wire [31:0] p2_smul_57594_comb;
  wire [31:0] p2_smul_57595_comb;
  wire [31:0] p2_smul_57596_comb;
  wire [31:0] p2_smul_57597_comb;
  wire [31:0] p2_smul_57598_comb;
  wire [31:0] p2_smul_57599_comb;
  wire [31:0] p2_smul_57600_comb;
  wire [31:0] p2_smul_57585_comb;
  wire [31:0] p2_smul_57586_comb;
  wire [31:0] p2_smul_57587_comb;
  wire [31:0] p2_smul_57588_comb;
  wire [31:0] p2_smul_57589_comb;
  wire [31:0] p2_smul_57590_comb;
  wire [31:0] p2_smul_57591_comb;
  wire [31:0] p2_smul_57592_comb;
  wire [31:0] p2_smul_57577_comb;
  wire [31:0] p2_smul_57578_comb;
  wire [31:0] p2_smul_57579_comb;
  wire [31:0] p2_smul_57580_comb;
  wire [31:0] p2_smul_57581_comb;
  wire [31:0] p2_smul_57582_comb;
  wire [31:0] p2_smul_57583_comb;
  wire [31:0] p2_smul_57584_comb;
  wire [31:0] p2_smul_57569_comb;
  wire [31:0] p2_smul_57570_comb;
  wire [31:0] p2_smul_57571_comb;
  wire [31:0] p2_smul_57572_comb;
  wire [31:0] p2_smul_57573_comb;
  wire [31:0] p2_smul_57574_comb;
  wire [31:0] p2_smul_57575_comb;
  wire [31:0] p2_smul_57576_comb;
  wire [31:0] p2_smul_57561_comb;
  wire [31:0] p2_smul_57562_comb;
  wire [31:0] p2_smul_57563_comb;
  wire [31:0] p2_smul_57564_comb;
  wire [31:0] p2_smul_57565_comb;
  wire [31:0] p2_smul_57566_comb;
  wire [31:0] p2_smul_57567_comb;
  wire [31:0] p2_smul_57568_comb;
  wire [31:0] p2_smul_57553_comb;
  wire [31:0] p2_smul_57554_comb;
  wire [31:0] p2_smul_57555_comb;
  wire [31:0] p2_smul_57556_comb;
  wire [31:0] p2_smul_57557_comb;
  wire [31:0] p2_smul_57558_comb;
  wire [31:0] p2_smul_57559_comb;
  wire [31:0] p2_smul_57560_comb;
  wire [31:0] p2_smul_57545_comb;
  wire [31:0] p2_smul_57546_comb;
  wire [31:0] p2_smul_57547_comb;
  wire [31:0] p2_smul_57548_comb;
  wire [31:0] p2_smul_57549_comb;
  wire [31:0] p2_smul_57550_comb;
  wire [31:0] p2_smul_57551_comb;
  wire [31:0] p2_smul_57552_comb;
  wire [31:0] p2_smul_57537_comb;
  wire [31:0] p2_smul_57538_comb;
  wire [31:0] p2_smul_57539_comb;
  wire [31:0] p2_smul_57540_comb;
  wire [31:0] p2_smul_57541_comb;
  wire [31:0] p2_smul_57542_comb;
  wire [31:0] p2_smul_57543_comb;
  wire [31:0] p2_smul_57544_comb;
  wire [31:0] p2_smul_57529_comb;
  wire [31:0] p2_smul_57530_comb;
  wire [31:0] p2_smul_57531_comb;
  wire [31:0] p2_smul_57532_comb;
  wire [31:0] p2_smul_57533_comb;
  wire [31:0] p2_smul_57534_comb;
  wire [31:0] p2_smul_57535_comb;
  wire [31:0] p2_smul_57536_comb;
  wire [31:0] p2_smul_57521_comb;
  wire [31:0] p2_smul_57522_comb;
  wire [31:0] p2_smul_57523_comb;
  wire [31:0] p2_smul_57524_comb;
  wire [31:0] p2_smul_57525_comb;
  wire [31:0] p2_smul_57526_comb;
  wire [31:0] p2_smul_57527_comb;
  wire [31:0] p2_smul_57528_comb;
  wire [31:0] p2_smul_57513_comb;
  wire [31:0] p2_smul_57514_comb;
  wire [31:0] p2_smul_57515_comb;
  wire [31:0] p2_smul_57516_comb;
  wire [31:0] p2_smul_57517_comb;
  wire [31:0] p2_smul_57518_comb;
  wire [31:0] p2_smul_57519_comb;
  wire [31:0] p2_smul_57520_comb;
  wire [31:0] p2_smul_57505_comb;
  wire [31:0] p2_smul_57506_comb;
  wire [31:0] p2_smul_57507_comb;
  wire [31:0] p2_smul_57508_comb;
  wire [31:0] p2_smul_57509_comb;
  wire [31:0] p2_smul_57510_comb;
  wire [31:0] p2_smul_57511_comb;
  wire [31:0] p2_smul_57512_comb;
  wire [31:0] p2_smul_57497_comb;
  wire [31:0] p2_smul_57498_comb;
  wire [31:0] p2_smul_57499_comb;
  wire [31:0] p2_smul_57500_comb;
  wire [31:0] p2_smul_57501_comb;
  wire [31:0] p2_smul_57502_comb;
  wire [31:0] p2_smul_57503_comb;
  wire [31:0] p2_smul_57504_comb;
  wire [31:0] p2_smul_57489_comb;
  wire [31:0] p2_smul_57490_comb;
  wire [31:0] p2_smul_57491_comb;
  wire [31:0] p2_smul_57492_comb;
  wire [31:0] p2_smul_57493_comb;
  wire [31:0] p2_smul_57494_comb;
  wire [31:0] p2_smul_57495_comb;
  wire [31:0] p2_smul_57496_comb;
  wire [31:0] p2_smul_57481_comb;
  wire [31:0] p2_smul_57482_comb;
  wire [31:0] p2_smul_57483_comb;
  wire [31:0] p2_smul_57484_comb;
  wire [31:0] p2_smul_57485_comb;
  wire [31:0] p2_smul_57486_comb;
  wire [31:0] p2_smul_57487_comb;
  wire [31:0] p2_smul_57488_comb;
  wire [31:0] p2_smul_57473_comb;
  wire [31:0] p2_smul_57474_comb;
  wire [31:0] p2_smul_57475_comb;
  wire [31:0] p2_smul_57476_comb;
  wire [31:0] p2_smul_57477_comb;
  wire [31:0] p2_smul_57478_comb;
  wire [31:0] p2_smul_57479_comb;
  wire [31:0] p2_smul_57480_comb;
  wire [31:0] p2_smul_57465_comb;
  wire [31:0] p2_smul_57466_comb;
  wire [31:0] p2_smul_57467_comb;
  wire [31:0] p2_smul_57468_comb;
  wire [31:0] p2_smul_57469_comb;
  wire [31:0] p2_smul_57470_comb;
  wire [31:0] p2_smul_57471_comb;
  wire [31:0] p2_smul_57472_comb;
  wire [31:0] p2_smul_57457_comb;
  wire [31:0] p2_smul_57458_comb;
  wire [31:0] p2_smul_57459_comb;
  wire [31:0] p2_smul_57460_comb;
  wire [31:0] p2_smul_57461_comb;
  wire [31:0] p2_smul_57462_comb;
  wire [31:0] p2_smul_57463_comb;
  wire [31:0] p2_smul_57464_comb;
  wire [31:0] p2_smul_57449_comb;
  wire [31:0] p2_smul_57450_comb;
  wire [31:0] p2_smul_57451_comb;
  wire [31:0] p2_smul_57452_comb;
  wire [31:0] p2_smul_57453_comb;
  wire [31:0] p2_smul_57454_comb;
  wire [31:0] p2_smul_57455_comb;
  wire [31:0] p2_smul_57456_comb;
  wire [31:0] p2_smul_57441_comb;
  wire [31:0] p2_smul_57442_comb;
  wire [31:0] p2_smul_57443_comb;
  wire [31:0] p2_smul_57444_comb;
  wire [31:0] p2_smul_57445_comb;
  wire [31:0] p2_smul_57446_comb;
  wire [31:0] p2_smul_57447_comb;
  wire [31:0] p2_smul_57448_comb;
  wire [31:0] p2_smul_57433_comb;
  wire [31:0] p2_smul_57434_comb;
  wire [31:0] p2_smul_57435_comb;
  wire [31:0] p2_smul_57436_comb;
  wire [31:0] p2_smul_57437_comb;
  wire [31:0] p2_smul_57438_comb;
  wire [31:0] p2_smul_57439_comb;
  wire [31:0] p2_smul_57440_comb;
  wire [31:0] p2_smul_57425_comb;
  wire [31:0] p2_smul_57426_comb;
  wire [31:0] p2_smul_57427_comb;
  wire [31:0] p2_smul_57428_comb;
  wire [31:0] p2_smul_57429_comb;
  wire [31:0] p2_smul_57430_comb;
  wire [31:0] p2_smul_57431_comb;
  wire [31:0] p2_smul_57432_comb;
  wire [31:0] p2_smul_57417_comb;
  wire [31:0] p2_smul_57418_comb;
  wire [31:0] p2_smul_57419_comb;
  wire [31:0] p2_smul_57420_comb;
  wire [31:0] p2_smul_57421_comb;
  wire [31:0] p2_smul_57422_comb;
  wire [31:0] p2_smul_57423_comb;
  wire [31:0] p2_smul_57424_comb;
  wire [31:0] p2_smul_57409_comb;
  wire [31:0] p2_smul_57410_comb;
  wire [31:0] p2_smul_57411_comb;
  wire [31:0] p2_smul_57412_comb;
  wire [31:0] p2_smul_57413_comb;
  wire [31:0] p2_smul_57414_comb;
  wire [31:0] p2_smul_57415_comb;
  wire [31:0] p2_smul_57416_comb;
  wire [31:0] p2_smul_57401_comb;
  wire [31:0] p2_smul_57402_comb;
  wire [31:0] p2_smul_57403_comb;
  wire [31:0] p2_smul_57404_comb;
  wire [31:0] p2_smul_57405_comb;
  wire [31:0] p2_smul_57406_comb;
  wire [31:0] p2_smul_57407_comb;
  wire [31:0] p2_smul_57408_comb;
  wire [31:0] p2_smul_57393_comb;
  wire [31:0] p2_smul_57394_comb;
  wire [31:0] p2_smul_57395_comb;
  wire [31:0] p2_smul_57396_comb;
  wire [31:0] p2_smul_57397_comb;
  wire [31:0] p2_smul_57398_comb;
  wire [31:0] p2_smul_57399_comb;
  wire [31:0] p2_smul_57400_comb;
  wire [31:0] p2_smul_57385_comb;
  wire [31:0] p2_smul_57386_comb;
  wire [31:0] p2_smul_57387_comb;
  wire [31:0] p2_smul_57388_comb;
  wire [31:0] p2_smul_57389_comb;
  wire [31:0] p2_smul_57390_comb;
  wire [31:0] p2_smul_57391_comb;
  wire [31:0] p2_smul_57392_comb;
  wire [31:0] p2_smul_57377_comb;
  wire [31:0] p2_smul_57378_comb;
  wire [31:0] p2_smul_57379_comb;
  wire [31:0] p2_smul_57380_comb;
  wire [31:0] p2_smul_57381_comb;
  wire [31:0] p2_smul_57382_comb;
  wire [31:0] p2_smul_57383_comb;
  wire [31:0] p2_smul_57384_comb;
  wire [31:0] p2_smul_57369_comb;
  wire [31:0] p2_smul_57370_comb;
  wire [31:0] p2_smul_57371_comb;
  wire [31:0] p2_smul_57372_comb;
  wire [31:0] p2_smul_57373_comb;
  wire [31:0] p2_smul_57374_comb;
  wire [31:0] p2_smul_57375_comb;
  wire [31:0] p2_smul_57376_comb;
  wire [31:0] p2_smul_57361_comb;
  wire [31:0] p2_smul_57362_comb;
  wire [31:0] p2_smul_57363_comb;
  wire [31:0] p2_smul_57364_comb;
  wire [31:0] p2_smul_57365_comb;
  wire [31:0] p2_smul_57366_comb;
  wire [31:0] p2_smul_57367_comb;
  wire [31:0] p2_smul_57368_comb;
  wire [31:0] p2_smul_57353_comb;
  wire [31:0] p2_smul_57354_comb;
  wire [31:0] p2_smul_57355_comb;
  wire [31:0] p2_smul_57356_comb;
  wire [31:0] p2_smul_57357_comb;
  wire [31:0] p2_smul_57358_comb;
  wire [31:0] p2_smul_57359_comb;
  wire [31:0] p2_smul_57360_comb;
  wire [31:0] p2_smul_57345_comb;
  wire [31:0] p2_smul_57346_comb;
  wire [31:0] p2_smul_57347_comb;
  wire [31:0] p2_smul_57348_comb;
  wire [31:0] p2_smul_57349_comb;
  wire [31:0] p2_smul_57350_comb;
  wire [31:0] p2_smul_57351_comb;
  wire [31:0] p2_smul_57352_comb;
  wire [31:0] p2_smul_57337_comb;
  wire [31:0] p2_smul_57338_comb;
  wire [31:0] p2_smul_57339_comb;
  wire [31:0] p2_smul_57340_comb;
  wire [31:0] p2_smul_57341_comb;
  wire [31:0] p2_smul_57342_comb;
  wire [31:0] p2_smul_57343_comb;
  wire [31:0] p2_smul_57344_comb;
  wire [31:0] p2_add_58101_comb;
  wire [31:0] p2_add_58102_comb;
  wire [31:0] p2_add_58103_comb;
  wire [31:0] p2_add_58104_comb;
  wire [31:0] p2_add_58097_comb;
  wire [31:0] p2_add_58098_comb;
  wire [31:0] p2_add_58099_comb;
  wire [31:0] p2_add_58100_comb;
  wire [31:0] p2_add_58093_comb;
  wire [31:0] p2_add_58094_comb;
  wire [31:0] p2_add_58095_comb;
  wire [31:0] p2_add_58096_comb;
  wire [31:0] p2_add_58089_comb;
  wire [31:0] p2_add_58090_comb;
  wire [31:0] p2_add_58091_comb;
  wire [31:0] p2_add_58092_comb;
  wire [31:0] p2_add_58085_comb;
  wire [31:0] p2_add_58086_comb;
  wire [31:0] p2_add_58087_comb;
  wire [31:0] p2_add_58088_comb;
  wire [31:0] p2_add_58081_comb;
  wire [31:0] p2_add_58082_comb;
  wire [31:0] p2_add_58083_comb;
  wire [31:0] p2_add_58084_comb;
  wire [31:0] p2_add_58077_comb;
  wire [31:0] p2_add_58078_comb;
  wire [31:0] p2_add_58079_comb;
  wire [31:0] p2_add_58080_comb;
  wire [31:0] p2_add_58073_comb;
  wire [31:0] p2_add_58074_comb;
  wire [31:0] p2_add_58075_comb;
  wire [31:0] p2_add_58076_comb;
  wire [31:0] p2_add_58069_comb;
  wire [31:0] p2_add_58070_comb;
  wire [31:0] p2_add_58071_comb;
  wire [31:0] p2_add_58072_comb;
  wire [31:0] p2_add_58065_comb;
  wire [31:0] p2_add_58066_comb;
  wire [31:0] p2_add_58067_comb;
  wire [31:0] p2_add_58068_comb;
  wire [31:0] p2_add_58061_comb;
  wire [31:0] p2_add_58062_comb;
  wire [31:0] p2_add_58063_comb;
  wire [31:0] p2_add_58064_comb;
  wire [31:0] p2_add_58057_comb;
  wire [31:0] p2_add_58058_comb;
  wire [31:0] p2_add_58059_comb;
  wire [31:0] p2_add_58060_comb;
  wire [31:0] p2_add_58053_comb;
  wire [31:0] p2_add_58054_comb;
  wire [31:0] p2_add_58055_comb;
  wire [31:0] p2_add_58056_comb;
  wire [31:0] p2_add_58049_comb;
  wire [31:0] p2_add_58050_comb;
  wire [31:0] p2_add_58051_comb;
  wire [31:0] p2_add_58052_comb;
  wire [31:0] p2_add_58045_comb;
  wire [31:0] p2_add_58046_comb;
  wire [31:0] p2_add_58047_comb;
  wire [31:0] p2_add_58048_comb;
  wire [31:0] p2_add_58041_comb;
  wire [31:0] p2_add_58042_comb;
  wire [31:0] p2_add_58043_comb;
  wire [31:0] p2_add_58044_comb;
  wire [31:0] p2_add_58037_comb;
  wire [31:0] p2_add_58038_comb;
  wire [31:0] p2_add_58039_comb;
  wire [31:0] p2_add_58040_comb;
  wire [31:0] p2_add_58033_comb;
  wire [31:0] p2_add_58034_comb;
  wire [31:0] p2_add_58035_comb;
  wire [31:0] p2_add_58036_comb;
  wire [31:0] p2_add_58029_comb;
  wire [31:0] p2_add_58030_comb;
  wire [31:0] p2_add_58031_comb;
  wire [31:0] p2_add_58032_comb;
  wire [31:0] p2_add_58025_comb;
  wire [31:0] p2_add_58026_comb;
  wire [31:0] p2_add_58027_comb;
  wire [31:0] p2_add_58028_comb;
  wire [31:0] p2_add_58021_comb;
  wire [31:0] p2_add_58022_comb;
  wire [31:0] p2_add_58023_comb;
  wire [31:0] p2_add_58024_comb;
  wire [31:0] p2_add_58017_comb;
  wire [31:0] p2_add_58018_comb;
  wire [31:0] p2_add_58019_comb;
  wire [31:0] p2_add_58020_comb;
  wire [31:0] p2_add_58013_comb;
  wire [31:0] p2_add_58014_comb;
  wire [31:0] p2_add_58015_comb;
  wire [31:0] p2_add_58016_comb;
  wire [31:0] p2_add_58009_comb;
  wire [31:0] p2_add_58010_comb;
  wire [31:0] p2_add_58011_comb;
  wire [31:0] p2_add_58012_comb;
  wire [31:0] p2_add_58005_comb;
  wire [31:0] p2_add_58006_comb;
  wire [31:0] p2_add_58007_comb;
  wire [31:0] p2_add_58008_comb;
  wire [31:0] p2_add_58001_comb;
  wire [31:0] p2_add_58002_comb;
  wire [31:0] p2_add_58003_comb;
  wire [31:0] p2_add_58004_comb;
  wire [31:0] p2_add_57997_comb;
  wire [31:0] p2_add_57998_comb;
  wire [31:0] p2_add_57999_comb;
  wire [31:0] p2_add_58000_comb;
  wire [31:0] p2_add_57993_comb;
  wire [31:0] p2_add_57994_comb;
  wire [31:0] p2_add_57995_comb;
  wire [31:0] p2_add_57996_comb;
  wire [31:0] p2_add_57989_comb;
  wire [31:0] p2_add_57990_comb;
  wire [31:0] p2_add_57991_comb;
  wire [31:0] p2_add_57992_comb;
  wire [31:0] p2_add_57985_comb;
  wire [31:0] p2_add_57986_comb;
  wire [31:0] p2_add_57987_comb;
  wire [31:0] p2_add_57988_comb;
  wire [31:0] p2_add_57981_comb;
  wire [31:0] p2_add_57982_comb;
  wire [31:0] p2_add_57983_comb;
  wire [31:0] p2_add_57984_comb;
  wire [31:0] p2_add_57977_comb;
  wire [31:0] p2_add_57978_comb;
  wire [31:0] p2_add_57979_comb;
  wire [31:0] p2_add_57980_comb;
  wire [31:0] p2_add_57973_comb;
  wire [31:0] p2_add_57974_comb;
  wire [31:0] p2_add_57975_comb;
  wire [31:0] p2_add_57976_comb;
  wire [31:0] p2_add_57969_comb;
  wire [31:0] p2_add_57970_comb;
  wire [31:0] p2_add_57971_comb;
  wire [31:0] p2_add_57972_comb;
  wire [31:0] p2_add_57965_comb;
  wire [31:0] p2_add_57966_comb;
  wire [31:0] p2_add_57967_comb;
  wire [31:0] p2_add_57968_comb;
  wire [31:0] p2_add_57961_comb;
  wire [31:0] p2_add_57962_comb;
  wire [31:0] p2_add_57963_comb;
  wire [31:0] p2_add_57964_comb;
  wire [31:0] p2_add_57957_comb;
  wire [31:0] p2_add_57958_comb;
  wire [31:0] p2_add_57959_comb;
  wire [31:0] p2_add_57960_comb;
  wire [31:0] p2_add_57953_comb;
  wire [31:0] p2_add_57954_comb;
  wire [31:0] p2_add_57955_comb;
  wire [31:0] p2_add_57956_comb;
  wire [31:0] p2_add_57949_comb;
  wire [31:0] p2_add_57950_comb;
  wire [31:0] p2_add_57951_comb;
  wire [31:0] p2_add_57952_comb;
  wire [31:0] p2_add_57945_comb;
  wire [31:0] p2_add_57946_comb;
  wire [31:0] p2_add_57947_comb;
  wire [31:0] p2_add_57948_comb;
  wire [31:0] p2_add_57941_comb;
  wire [31:0] p2_add_57942_comb;
  wire [31:0] p2_add_57943_comb;
  wire [31:0] p2_add_57944_comb;
  wire [31:0] p2_add_57937_comb;
  wire [31:0] p2_add_57938_comb;
  wire [31:0] p2_add_57939_comb;
  wire [31:0] p2_add_57940_comb;
  wire [31:0] p2_add_57933_comb;
  wire [31:0] p2_add_57934_comb;
  wire [31:0] p2_add_57935_comb;
  wire [31:0] p2_add_57936_comb;
  wire [31:0] p2_add_57929_comb;
  wire [31:0] p2_add_57930_comb;
  wire [31:0] p2_add_57931_comb;
  wire [31:0] p2_add_57932_comb;
  wire [31:0] p2_add_57925_comb;
  wire [31:0] p2_add_57926_comb;
  wire [31:0] p2_add_57927_comb;
  wire [31:0] p2_add_57928_comb;
  wire [31:0] p2_add_57921_comb;
  wire [31:0] p2_add_57922_comb;
  wire [31:0] p2_add_57923_comb;
  wire [31:0] p2_add_57924_comb;
  wire [31:0] p2_add_57917_comb;
  wire [31:0] p2_add_57918_comb;
  wire [31:0] p2_add_57919_comb;
  wire [31:0] p2_add_57920_comb;
  wire [31:0] p2_add_57913_comb;
  wire [31:0] p2_add_57914_comb;
  wire [31:0] p2_add_57915_comb;
  wire [31:0] p2_add_57916_comb;
  wire [31:0] p2_add_57909_comb;
  wire [31:0] p2_add_57910_comb;
  wire [31:0] p2_add_57911_comb;
  wire [31:0] p2_add_57912_comb;
  wire [31:0] p2_add_57905_comb;
  wire [31:0] p2_add_57906_comb;
  wire [31:0] p2_add_57907_comb;
  wire [31:0] p2_add_57908_comb;
  wire [31:0] p2_add_57901_comb;
  wire [31:0] p2_add_57902_comb;
  wire [31:0] p2_add_57903_comb;
  wire [31:0] p2_add_57904_comb;
  wire [31:0] p2_add_57897_comb;
  wire [31:0] p2_add_57898_comb;
  wire [31:0] p2_add_57899_comb;
  wire [31:0] p2_add_57900_comb;
  wire [31:0] p2_add_57893_comb;
  wire [31:0] p2_add_57894_comb;
  wire [31:0] p2_add_57895_comb;
  wire [31:0] p2_add_57896_comb;
  wire [31:0] p2_add_57889_comb;
  wire [31:0] p2_add_57890_comb;
  wire [31:0] p2_add_57891_comb;
  wire [31:0] p2_add_57892_comb;
  wire [31:0] p2_add_57885_comb;
  wire [31:0] p2_add_57886_comb;
  wire [31:0] p2_add_57887_comb;
  wire [31:0] p2_add_57888_comb;
  wire [31:0] p2_add_57881_comb;
  wire [31:0] p2_add_57882_comb;
  wire [31:0] p2_add_57883_comb;
  wire [31:0] p2_add_57884_comb;
  wire [31:0] p2_add_57877_comb;
  wire [31:0] p2_add_57878_comb;
  wire [31:0] p2_add_57879_comb;
  wire [31:0] p2_add_57880_comb;
  wire [31:0] p2_add_57873_comb;
  wire [31:0] p2_add_57874_comb;
  wire [31:0] p2_add_57875_comb;
  wire [31:0] p2_add_57876_comb;
  wire [31:0] p2_add_57869_comb;
  wire [31:0] p2_add_57870_comb;
  wire [31:0] p2_add_57871_comb;
  wire [31:0] p2_add_57872_comb;
  wire [31:0] p2_add_57865_comb;
  wire [31:0] p2_add_57866_comb;
  wire [31:0] p2_add_57867_comb;
  wire [31:0] p2_add_57868_comb;
  wire [31:0] p2_add_57861_comb;
  wire [31:0] p2_add_57862_comb;
  wire [31:0] p2_add_57863_comb;
  wire [31:0] p2_add_57864_comb;
  wire [31:0] p2_add_57857_comb;
  wire [31:0] p2_add_57858_comb;
  wire [31:0] p2_add_57859_comb;
  wire [31:0] p2_add_57860_comb;
  wire [31:0] p2_add_57853_comb;
  wire [31:0] p2_add_57854_comb;
  wire [31:0] p2_add_57855_comb;
  wire [31:0] p2_add_57856_comb;
  wire [31:0] p2_add_57849_comb;
  wire [31:0] p2_add_57850_comb;
  wire [31:0] p2_add_57851_comb;
  wire [31:0] p2_add_57852_comb;
  assign p2_smul_57841_comb = smul32b_32b_x_32b(p1_array_index_57069, p1_array_index_57013);
  assign p2_smul_57842_comb = smul32b_32b_x_32b(p1_array_index_57070, p1_array_index_57014);
  assign p2_smul_57843_comb = smul32b_32b_x_32b(p1_array_index_57071, p1_array_index_57015);
  assign p2_smul_57844_comb = smul32b_32b_x_32b(p1_array_index_57072, p1_array_index_57016);
  assign p2_smul_57845_comb = smul32b_32b_x_32b(p1_array_index_57076, p1_array_index_57017);
  assign p2_smul_57846_comb = smul32b_32b_x_32b(p1_array_index_57075, p1_array_index_57018);
  assign p2_smul_57847_comb = smul32b_32b_x_32b(p1_array_index_57074, p1_array_index_57019);
  assign p2_smul_57848_comb = smul32b_32b_x_32b(p1_array_index_57073, p1_array_index_57020);
  assign p2_smul_57833_comb = smul32b_32b_x_32b(p1_array_index_57069, p1_array_index_57005);
  assign p2_smul_57834_comb = smul32b_32b_x_32b(p1_array_index_57070, p1_array_index_57006);
  assign p2_smul_57835_comb = smul32b_32b_x_32b(p1_array_index_57071, p1_array_index_57007);
  assign p2_smul_57836_comb = smul32b_32b_x_32b(p1_array_index_57072, p1_array_index_57008);
  assign p2_smul_57837_comb = smul32b_32b_x_32b(p1_array_index_57076, p1_array_index_57012);
  assign p2_smul_57838_comb = smul32b_32b_x_32b(p1_array_index_57075, p1_array_index_57011);
  assign p2_smul_57839_comb = smul32b_32b_x_32b(p1_array_index_57074, p1_array_index_57010);
  assign p2_smul_57840_comb = smul32b_32b_x_32b(p1_array_index_57073, p1_array_index_57009);
  assign p2_smul_57825_comb = smul32b_32b_x_32b(p1_array_index_57069, p1_array_index_56997);
  assign p2_smul_57826_comb = smul32b_32b_x_32b(p1_array_index_57070, p1_array_index_56998);
  assign p2_smul_57827_comb = smul32b_32b_x_32b(p1_array_index_57071, p1_array_index_56999);
  assign p2_smul_57828_comb = smul32b_32b_x_32b(p1_array_index_57072, p1_array_index_57000);
  assign p2_smul_57829_comb = smul32b_32b_x_32b(p1_array_index_57076, p1_array_index_57001);
  assign p2_smul_57830_comb = smul32b_32b_x_32b(p1_array_index_57075, p1_array_index_57002);
  assign p2_smul_57831_comb = smul32b_32b_x_32b(p1_array_index_57074, p1_array_index_57003);
  assign p2_smul_57832_comb = smul32b_32b_x_32b(p1_array_index_57073, p1_array_index_57004);
  assign p2_smul_57817_comb = smul32b_32b_x_32b(p1_array_index_57069, p1_array_index_56989);
  assign p2_smul_57818_comb = smul32b_32b_x_32b(p1_array_index_57070, p1_array_index_56990);
  assign p2_smul_57819_comb = smul32b_32b_x_32b(p1_array_index_57071, p1_array_index_56991);
  assign p2_smul_57820_comb = smul32b_32b_x_32b(p1_array_index_57072, p1_array_index_56992);
  assign p2_smul_57821_comb = smul32b_32b_x_32b(p1_array_index_57076, p1_array_index_56993);
  assign p2_smul_57822_comb = smul32b_32b_x_32b(p1_array_index_57075, p1_array_index_56994);
  assign p2_smul_57823_comb = smul32b_32b_x_32b(p1_array_index_57074, p1_array_index_56995);
  assign p2_smul_57824_comb = smul32b_32b_x_32b(p1_array_index_57073, p1_array_index_56996);
  assign p2_smul_57809_comb = smul32b_32b_x_32b(p1_array_index_57069, p1_array_index_56981);
  assign p2_smul_57810_comb = smul32b_32b_x_32b(p1_array_index_57070, p1_array_index_56982);
  assign p2_smul_57811_comb = smul32b_32b_x_32b(p1_array_index_57071, p1_array_index_56983);
  assign p2_smul_57812_comb = smul32b_32b_x_32b(p1_array_index_57072, p1_array_index_56984);
  assign p2_smul_57813_comb = smul32b_32b_x_32b(p1_array_index_57076, p1_array_index_56985);
  assign p2_smul_57814_comb = smul32b_32b_x_32b(p1_array_index_57075, p1_array_index_56986);
  assign p2_smul_57815_comb = smul32b_32b_x_32b(p1_array_index_57074, p1_array_index_56987);
  assign p2_smul_57816_comb = smul32b_32b_x_32b(p1_array_index_57073, p1_array_index_56988);
  assign p2_smul_57801_comb = smul32b_32b_x_32b(p1_array_index_57069, p1_array_index_56973);
  assign p2_smul_57802_comb = smul32b_32b_x_32b(p1_array_index_57070, p1_array_index_56974);
  assign p2_smul_57803_comb = smul32b_32b_x_32b(p1_array_index_57071, p1_array_index_56975);
  assign p2_smul_57804_comb = smul32b_32b_x_32b(p1_array_index_57072, p1_array_index_56976);
  assign p2_smul_57805_comb = smul32b_32b_x_32b(p1_array_index_57076, p1_array_index_56977);
  assign p2_smul_57806_comb = smul32b_32b_x_32b(p1_array_index_57075, p1_array_index_56978);
  assign p2_smul_57807_comb = smul32b_32b_x_32b(p1_array_index_57074, p1_array_index_56979);
  assign p2_smul_57808_comb = smul32b_32b_x_32b(p1_array_index_57073, p1_array_index_56980);
  assign p2_smul_57793_comb = smul32b_32b_x_32b(p1_array_index_57069, p1_array_index_56965);
  assign p2_smul_57794_comb = smul32b_32b_x_32b(p1_array_index_57070, p1_array_index_56966);
  assign p2_smul_57795_comb = smul32b_32b_x_32b(p1_array_index_57071, p1_array_index_56967);
  assign p2_smul_57796_comb = smul32b_32b_x_32b(p1_array_index_57072, p1_array_index_56968);
  assign p2_smul_57797_comb = smul32b_32b_x_32b(p1_array_index_57076, p1_array_index_56969);
  assign p2_smul_57798_comb = smul32b_32b_x_32b(p1_array_index_57075, p1_array_index_56970);
  assign p2_smul_57799_comb = smul32b_32b_x_32b(p1_array_index_57074, p1_array_index_56971);
  assign p2_smul_57800_comb = smul32b_32b_x_32b(p1_array_index_57073, p1_array_index_56972);
  assign p2_smul_57785_comb = smul32b_32b_x_32b(p1_array_index_57069, p1_array_index_56950);
  assign p2_smul_57786_comb = smul32b_32b_x_32b(p1_array_index_57070, p1_array_index_56952);
  assign p2_smul_57787_comb = smul32b_32b_x_32b(p1_array_index_57071, p1_array_index_56954);
  assign p2_smul_57788_comb = smul32b_32b_x_32b(p1_array_index_57072, p1_array_index_56956);
  assign p2_smul_57789_comb = smul32b_32b_x_32b(p1_array_index_57073, p1_array_index_56964);
  assign p2_smul_57790_comb = smul32b_32b_x_32b(p1_array_index_57074, p1_array_index_56962);
  assign p2_smul_57791_comb = smul32b_32b_x_32b(p1_array_index_57075, p1_array_index_56960);
  assign p2_smul_57792_comb = smul32b_32b_x_32b(p1_array_index_57076, p1_array_index_56958);
  assign p2_smul_57777_comb = smul32b_32b_x_32b(p1_array_index_57061, p1_array_index_57013);
  assign p2_smul_57778_comb = smul32b_32b_x_32b(p1_array_index_57062, p1_array_index_57014);
  assign p2_smul_57779_comb = smul32b_32b_x_32b(p1_array_index_57063, p1_array_index_57015);
  assign p2_smul_57780_comb = smul32b_32b_x_32b(p1_array_index_57064, p1_array_index_57016);
  assign p2_smul_57781_comb = smul32b_32b_x_32b(p1_array_index_57065, p1_array_index_57017);
  assign p2_smul_57782_comb = smul32b_32b_x_32b(p1_array_index_57066, p1_array_index_57018);
  assign p2_smul_57783_comb = smul32b_32b_x_32b(p1_array_index_57067, p1_array_index_57019);
  assign p2_smul_57784_comb = smul32b_32b_x_32b(p1_array_index_57068, p1_array_index_57020);
  assign p2_smul_57769_comb = smul32b_32b_x_32b(p1_array_index_57061, p1_array_index_57005);
  assign p2_smul_57770_comb = smul32b_32b_x_32b(p1_array_index_57062, p1_array_index_57006);
  assign p2_smul_57771_comb = smul32b_32b_x_32b(p1_array_index_57063, p1_array_index_57007);
  assign p2_smul_57772_comb = smul32b_32b_x_32b(p1_array_index_57064, p1_array_index_57008);
  assign p2_smul_57773_comb = smul32b_32b_x_32b(p1_array_index_57065, p1_array_index_57012);
  assign p2_smul_57774_comb = smul32b_32b_x_32b(p1_array_index_57066, p1_array_index_57011);
  assign p2_smul_57775_comb = smul32b_32b_x_32b(p1_array_index_57067, p1_array_index_57010);
  assign p2_smul_57776_comb = smul32b_32b_x_32b(p1_array_index_57068, p1_array_index_57009);
  assign p2_smul_57761_comb = smul32b_32b_x_32b(p1_array_index_57061, p1_array_index_56997);
  assign p2_smul_57762_comb = smul32b_32b_x_32b(p1_array_index_57062, p1_array_index_56998);
  assign p2_smul_57763_comb = smul32b_32b_x_32b(p1_array_index_57063, p1_array_index_56999);
  assign p2_smul_57764_comb = smul32b_32b_x_32b(p1_array_index_57064, p1_array_index_57000);
  assign p2_smul_57765_comb = smul32b_32b_x_32b(p1_array_index_57065, p1_array_index_57001);
  assign p2_smul_57766_comb = smul32b_32b_x_32b(p1_array_index_57066, p1_array_index_57002);
  assign p2_smul_57767_comb = smul32b_32b_x_32b(p1_array_index_57067, p1_array_index_57003);
  assign p2_smul_57768_comb = smul32b_32b_x_32b(p1_array_index_57068, p1_array_index_57004);
  assign p2_smul_57753_comb = smul32b_32b_x_32b(p1_array_index_57061, p1_array_index_56989);
  assign p2_smul_57754_comb = smul32b_32b_x_32b(p1_array_index_57062, p1_array_index_56990);
  assign p2_smul_57755_comb = smul32b_32b_x_32b(p1_array_index_57063, p1_array_index_56991);
  assign p2_smul_57756_comb = smul32b_32b_x_32b(p1_array_index_57064, p1_array_index_56992);
  assign p2_smul_57757_comb = smul32b_32b_x_32b(p1_array_index_57065, p1_array_index_56993);
  assign p2_smul_57758_comb = smul32b_32b_x_32b(p1_array_index_57066, p1_array_index_56994);
  assign p2_smul_57759_comb = smul32b_32b_x_32b(p1_array_index_57067, p1_array_index_56995);
  assign p2_smul_57760_comb = smul32b_32b_x_32b(p1_array_index_57068, p1_array_index_56996);
  assign p2_smul_57745_comb = smul32b_32b_x_32b(p1_array_index_57061, p1_array_index_56981);
  assign p2_smul_57746_comb = smul32b_32b_x_32b(p1_array_index_57062, p1_array_index_56982);
  assign p2_smul_57747_comb = smul32b_32b_x_32b(p1_array_index_57063, p1_array_index_56983);
  assign p2_smul_57748_comb = smul32b_32b_x_32b(p1_array_index_57064, p1_array_index_56984);
  assign p2_smul_57749_comb = smul32b_32b_x_32b(p1_array_index_57065, p1_array_index_56985);
  assign p2_smul_57750_comb = smul32b_32b_x_32b(p1_array_index_57066, p1_array_index_56986);
  assign p2_smul_57751_comb = smul32b_32b_x_32b(p1_array_index_57067, p1_array_index_56987);
  assign p2_smul_57752_comb = smul32b_32b_x_32b(p1_array_index_57068, p1_array_index_56988);
  assign p2_smul_57737_comb = smul32b_32b_x_32b(p1_array_index_57061, p1_array_index_56973);
  assign p2_smul_57738_comb = smul32b_32b_x_32b(p1_array_index_57062, p1_array_index_56974);
  assign p2_smul_57739_comb = smul32b_32b_x_32b(p1_array_index_57063, p1_array_index_56975);
  assign p2_smul_57740_comb = smul32b_32b_x_32b(p1_array_index_57064, p1_array_index_56976);
  assign p2_smul_57741_comb = smul32b_32b_x_32b(p1_array_index_57065, p1_array_index_56977);
  assign p2_smul_57742_comb = smul32b_32b_x_32b(p1_array_index_57066, p1_array_index_56978);
  assign p2_smul_57743_comb = smul32b_32b_x_32b(p1_array_index_57067, p1_array_index_56979);
  assign p2_smul_57744_comb = smul32b_32b_x_32b(p1_array_index_57068, p1_array_index_56980);
  assign p2_smul_57729_comb = smul32b_32b_x_32b(p1_array_index_57061, p1_array_index_56965);
  assign p2_smul_57730_comb = smul32b_32b_x_32b(p1_array_index_57062, p1_array_index_56966);
  assign p2_smul_57731_comb = smul32b_32b_x_32b(p1_array_index_57063, p1_array_index_56967);
  assign p2_smul_57732_comb = smul32b_32b_x_32b(p1_array_index_57064, p1_array_index_56968);
  assign p2_smul_57733_comb = smul32b_32b_x_32b(p1_array_index_57065, p1_array_index_56969);
  assign p2_smul_57734_comb = smul32b_32b_x_32b(p1_array_index_57066, p1_array_index_56970);
  assign p2_smul_57735_comb = smul32b_32b_x_32b(p1_array_index_57067, p1_array_index_56971);
  assign p2_smul_57736_comb = smul32b_32b_x_32b(p1_array_index_57068, p1_array_index_56972);
  assign p2_smul_57721_comb = smul32b_32b_x_32b(p1_array_index_57061, p1_array_index_56950);
  assign p2_smul_57722_comb = smul32b_32b_x_32b(p1_array_index_57062, p1_array_index_56952);
  assign p2_smul_57723_comb = smul32b_32b_x_32b(p1_array_index_57063, p1_array_index_56954);
  assign p2_smul_57724_comb = smul32b_32b_x_32b(p1_array_index_57064, p1_array_index_56956);
  assign p2_smul_57725_comb = smul32b_32b_x_32b(p1_array_index_57065, p1_array_index_56958);
  assign p2_smul_57726_comb = smul32b_32b_x_32b(p1_array_index_57066, p1_array_index_56960);
  assign p2_smul_57727_comb = smul32b_32b_x_32b(p1_array_index_57067, p1_array_index_56962);
  assign p2_smul_57728_comb = smul32b_32b_x_32b(p1_array_index_57068, p1_array_index_56964);
  assign p2_smul_57713_comb = smul32b_32b_x_32b(p1_array_index_57053, p1_array_index_57013);
  assign p2_smul_57714_comb = smul32b_32b_x_32b(p1_array_index_57054, p1_array_index_57014);
  assign p2_smul_57715_comb = smul32b_32b_x_32b(p1_array_index_57055, p1_array_index_57015);
  assign p2_smul_57716_comb = smul32b_32b_x_32b(p1_array_index_57056, p1_array_index_57016);
  assign p2_smul_57717_comb = smul32b_32b_x_32b(p1_array_index_57057, p1_array_index_57017);
  assign p2_smul_57718_comb = smul32b_32b_x_32b(p1_array_index_57058, p1_array_index_57018);
  assign p2_smul_57719_comb = smul32b_32b_x_32b(p1_array_index_57059, p1_array_index_57019);
  assign p2_smul_57720_comb = smul32b_32b_x_32b(p1_array_index_57060, p1_array_index_57020);
  assign p2_smul_57705_comb = smul32b_32b_x_32b(p1_array_index_57053, p1_array_index_57005);
  assign p2_smul_57706_comb = smul32b_32b_x_32b(p1_array_index_57054, p1_array_index_57006);
  assign p2_smul_57707_comb = smul32b_32b_x_32b(p1_array_index_57055, p1_array_index_57007);
  assign p2_smul_57708_comb = smul32b_32b_x_32b(p1_array_index_57056, p1_array_index_57008);
  assign p2_smul_57709_comb = smul32b_32b_x_32b(p1_array_index_57057, p1_array_index_57012);
  assign p2_smul_57710_comb = smul32b_32b_x_32b(p1_array_index_57058, p1_array_index_57011);
  assign p2_smul_57711_comb = smul32b_32b_x_32b(p1_array_index_57059, p1_array_index_57010);
  assign p2_smul_57712_comb = smul32b_32b_x_32b(p1_array_index_57060, p1_array_index_57009);
  assign p2_smul_57697_comb = smul32b_32b_x_32b(p1_array_index_57053, p1_array_index_56997);
  assign p2_smul_57698_comb = smul32b_32b_x_32b(p1_array_index_57054, p1_array_index_56998);
  assign p2_smul_57699_comb = smul32b_32b_x_32b(p1_array_index_57055, p1_array_index_56999);
  assign p2_smul_57700_comb = smul32b_32b_x_32b(p1_array_index_57056, p1_array_index_57000);
  assign p2_smul_57701_comb = smul32b_32b_x_32b(p1_array_index_57057, p1_array_index_57001);
  assign p2_smul_57702_comb = smul32b_32b_x_32b(p1_array_index_57058, p1_array_index_57002);
  assign p2_smul_57703_comb = smul32b_32b_x_32b(p1_array_index_57059, p1_array_index_57003);
  assign p2_smul_57704_comb = smul32b_32b_x_32b(p1_array_index_57060, p1_array_index_57004);
  assign p2_smul_57689_comb = smul32b_32b_x_32b(p1_array_index_57053, p1_array_index_56989);
  assign p2_smul_57690_comb = smul32b_32b_x_32b(p1_array_index_57054, p1_array_index_56990);
  assign p2_smul_57691_comb = smul32b_32b_x_32b(p1_array_index_57055, p1_array_index_56991);
  assign p2_smul_57692_comb = smul32b_32b_x_32b(p1_array_index_57056, p1_array_index_56992);
  assign p2_smul_57693_comb = smul32b_32b_x_32b(p1_array_index_57057, p1_array_index_56993);
  assign p2_smul_57694_comb = smul32b_32b_x_32b(p1_array_index_57058, p1_array_index_56994);
  assign p2_smul_57695_comb = smul32b_32b_x_32b(p1_array_index_57059, p1_array_index_56995);
  assign p2_smul_57696_comb = smul32b_32b_x_32b(p1_array_index_57060, p1_array_index_56996);
  assign p2_smul_57681_comb = smul32b_32b_x_32b(p1_array_index_57053, p1_array_index_56981);
  assign p2_smul_57682_comb = smul32b_32b_x_32b(p1_array_index_57054, p1_array_index_56982);
  assign p2_smul_57683_comb = smul32b_32b_x_32b(p1_array_index_57055, p1_array_index_56983);
  assign p2_smul_57684_comb = smul32b_32b_x_32b(p1_array_index_57056, p1_array_index_56984);
  assign p2_smul_57685_comb = smul32b_32b_x_32b(p1_array_index_57057, p1_array_index_56985);
  assign p2_smul_57686_comb = smul32b_32b_x_32b(p1_array_index_57058, p1_array_index_56986);
  assign p2_smul_57687_comb = smul32b_32b_x_32b(p1_array_index_57059, p1_array_index_56987);
  assign p2_smul_57688_comb = smul32b_32b_x_32b(p1_array_index_57060, p1_array_index_56988);
  assign p2_smul_57673_comb = smul32b_32b_x_32b(p1_array_index_57053, p1_array_index_56973);
  assign p2_smul_57674_comb = smul32b_32b_x_32b(p1_array_index_57054, p1_array_index_56974);
  assign p2_smul_57675_comb = smul32b_32b_x_32b(p1_array_index_57055, p1_array_index_56975);
  assign p2_smul_57676_comb = smul32b_32b_x_32b(p1_array_index_57056, p1_array_index_56976);
  assign p2_smul_57677_comb = smul32b_32b_x_32b(p1_array_index_57057, p1_array_index_56977);
  assign p2_smul_57678_comb = smul32b_32b_x_32b(p1_array_index_57058, p1_array_index_56978);
  assign p2_smul_57679_comb = smul32b_32b_x_32b(p1_array_index_57059, p1_array_index_56979);
  assign p2_smul_57680_comb = smul32b_32b_x_32b(p1_array_index_57060, p1_array_index_56980);
  assign p2_smul_57665_comb = smul32b_32b_x_32b(p1_array_index_57053, p1_array_index_56965);
  assign p2_smul_57666_comb = smul32b_32b_x_32b(p1_array_index_57054, p1_array_index_56966);
  assign p2_smul_57667_comb = smul32b_32b_x_32b(p1_array_index_57055, p1_array_index_56967);
  assign p2_smul_57668_comb = smul32b_32b_x_32b(p1_array_index_57056, p1_array_index_56968);
  assign p2_smul_57669_comb = smul32b_32b_x_32b(p1_array_index_57057, p1_array_index_56969);
  assign p2_smul_57670_comb = smul32b_32b_x_32b(p1_array_index_57058, p1_array_index_56970);
  assign p2_smul_57671_comb = smul32b_32b_x_32b(p1_array_index_57059, p1_array_index_56971);
  assign p2_smul_57672_comb = smul32b_32b_x_32b(p1_array_index_57060, p1_array_index_56972);
  assign p2_smul_57657_comb = smul32b_32b_x_32b(p1_array_index_57053, p1_array_index_56950);
  assign p2_smul_57658_comb = smul32b_32b_x_32b(p1_array_index_57054, p1_array_index_56952);
  assign p2_smul_57659_comb = smul32b_32b_x_32b(p1_array_index_57055, p1_array_index_56954);
  assign p2_smul_57660_comb = smul32b_32b_x_32b(p1_array_index_57056, p1_array_index_56956);
  assign p2_smul_57661_comb = smul32b_32b_x_32b(p1_array_index_57057, p1_array_index_56958);
  assign p2_smul_57662_comb = smul32b_32b_x_32b(p1_array_index_57058, p1_array_index_56960);
  assign p2_smul_57663_comb = smul32b_32b_x_32b(p1_array_index_57059, p1_array_index_56962);
  assign p2_smul_57664_comb = smul32b_32b_x_32b(p1_array_index_57060, p1_array_index_56964);
  assign p2_smul_57649_comb = smul32b_32b_x_32b(p1_array_index_57045, p1_array_index_57013);
  assign p2_smul_57650_comb = smul32b_32b_x_32b(p1_array_index_57046, p1_array_index_57014);
  assign p2_smul_57651_comb = smul32b_32b_x_32b(p1_array_index_57047, p1_array_index_57015);
  assign p2_smul_57652_comb = smul32b_32b_x_32b(p1_array_index_57048, p1_array_index_57016);
  assign p2_smul_57653_comb = smul32b_32b_x_32b(p1_array_index_57052, p1_array_index_57017);
  assign p2_smul_57654_comb = smul32b_32b_x_32b(p1_array_index_57051, p1_array_index_57018);
  assign p2_smul_57655_comb = smul32b_32b_x_32b(p1_array_index_57050, p1_array_index_57019);
  assign p2_smul_57656_comb = smul32b_32b_x_32b(p1_array_index_57049, p1_array_index_57020);
  assign p2_smul_57641_comb = smul32b_32b_x_32b(p1_array_index_57045, p1_array_index_57005);
  assign p2_smul_57642_comb = smul32b_32b_x_32b(p1_array_index_57046, p1_array_index_57006);
  assign p2_smul_57643_comb = smul32b_32b_x_32b(p1_array_index_57047, p1_array_index_57007);
  assign p2_smul_57644_comb = smul32b_32b_x_32b(p1_array_index_57048, p1_array_index_57008);
  assign p2_smul_57645_comb = smul32b_32b_x_32b(p1_array_index_57052, p1_array_index_57012);
  assign p2_smul_57646_comb = smul32b_32b_x_32b(p1_array_index_57051, p1_array_index_57011);
  assign p2_smul_57647_comb = smul32b_32b_x_32b(p1_array_index_57050, p1_array_index_57010);
  assign p2_smul_57648_comb = smul32b_32b_x_32b(p1_array_index_57049, p1_array_index_57009);
  assign p2_smul_57633_comb = smul32b_32b_x_32b(p1_array_index_57045, p1_array_index_56997);
  assign p2_smul_57634_comb = smul32b_32b_x_32b(p1_array_index_57046, p1_array_index_56998);
  assign p2_smul_57635_comb = smul32b_32b_x_32b(p1_array_index_57047, p1_array_index_56999);
  assign p2_smul_57636_comb = smul32b_32b_x_32b(p1_array_index_57048, p1_array_index_57000);
  assign p2_smul_57637_comb = smul32b_32b_x_32b(p1_array_index_57052, p1_array_index_57001);
  assign p2_smul_57638_comb = smul32b_32b_x_32b(p1_array_index_57051, p1_array_index_57002);
  assign p2_smul_57639_comb = smul32b_32b_x_32b(p1_array_index_57050, p1_array_index_57003);
  assign p2_smul_57640_comb = smul32b_32b_x_32b(p1_array_index_57049, p1_array_index_57004);
  assign p2_smul_57625_comb = smul32b_32b_x_32b(p1_array_index_57045, p1_array_index_56989);
  assign p2_smul_57626_comb = smul32b_32b_x_32b(p1_array_index_57046, p1_array_index_56990);
  assign p2_smul_57627_comb = smul32b_32b_x_32b(p1_array_index_57047, p1_array_index_56991);
  assign p2_smul_57628_comb = smul32b_32b_x_32b(p1_array_index_57048, p1_array_index_56992);
  assign p2_smul_57629_comb = smul32b_32b_x_32b(p1_array_index_57049, p1_array_index_56996);
  assign p2_smul_57630_comb = smul32b_32b_x_32b(p1_array_index_57050, p1_array_index_56995);
  assign p2_smul_57631_comb = smul32b_32b_x_32b(p1_array_index_57051, p1_array_index_56994);
  assign p2_smul_57632_comb = smul32b_32b_x_32b(p1_array_index_57052, p1_array_index_56993);
  assign p2_smul_57617_comb = smul32b_32b_x_32b(p1_array_index_57045, p1_array_index_56981);
  assign p2_smul_57618_comb = smul32b_32b_x_32b(p1_array_index_57046, p1_array_index_56982);
  assign p2_smul_57619_comb = smul32b_32b_x_32b(p1_array_index_57047, p1_array_index_56983);
  assign p2_smul_57620_comb = smul32b_32b_x_32b(p1_array_index_57048, p1_array_index_56984);
  assign p2_smul_57621_comb = smul32b_32b_x_32b(p1_array_index_57052, p1_array_index_56985);
  assign p2_smul_57622_comb = smul32b_32b_x_32b(p1_array_index_57051, p1_array_index_56986);
  assign p2_smul_57623_comb = smul32b_32b_x_32b(p1_array_index_57050, p1_array_index_56987);
  assign p2_smul_57624_comb = smul32b_32b_x_32b(p1_array_index_57049, p1_array_index_56988);
  assign p2_smul_57609_comb = smul32b_32b_x_32b(p1_array_index_57045, p1_array_index_56973);
  assign p2_smul_57610_comb = smul32b_32b_x_32b(p1_array_index_57046, p1_array_index_56974);
  assign p2_smul_57611_comb = smul32b_32b_x_32b(p1_array_index_57047, p1_array_index_56975);
  assign p2_smul_57612_comb = smul32b_32b_x_32b(p1_array_index_57048, p1_array_index_56976);
  assign p2_smul_57613_comb = smul32b_32b_x_32b(p1_array_index_57052, p1_array_index_56977);
  assign p2_smul_57614_comb = smul32b_32b_x_32b(p1_array_index_57051, p1_array_index_56978);
  assign p2_smul_57615_comb = smul32b_32b_x_32b(p1_array_index_57050, p1_array_index_56979);
  assign p2_smul_57616_comb = smul32b_32b_x_32b(p1_array_index_57049, p1_array_index_56980);
  assign p2_smul_57601_comb = smul32b_32b_x_32b(p1_array_index_57045, p1_array_index_56965);
  assign p2_smul_57602_comb = smul32b_32b_x_32b(p1_array_index_57046, p1_array_index_56966);
  assign p2_smul_57603_comb = smul32b_32b_x_32b(p1_array_index_57047, p1_array_index_56967);
  assign p2_smul_57604_comb = smul32b_32b_x_32b(p1_array_index_57048, p1_array_index_56968);
  assign p2_smul_57605_comb = smul32b_32b_x_32b(p1_array_index_57052, p1_array_index_56969);
  assign p2_smul_57606_comb = smul32b_32b_x_32b(p1_array_index_57051, p1_array_index_56970);
  assign p2_smul_57607_comb = smul32b_32b_x_32b(p1_array_index_57050, p1_array_index_56971);
  assign p2_smul_57608_comb = smul32b_32b_x_32b(p1_array_index_57049, p1_array_index_56972);
  assign p2_smul_57593_comb = smul32b_32b_x_32b(p1_array_index_57045, p1_array_index_56950);
  assign p2_smul_57594_comb = smul32b_32b_x_32b(p1_array_index_57046, p1_array_index_56952);
  assign p2_smul_57595_comb = smul32b_32b_x_32b(p1_array_index_57047, p1_array_index_56954);
  assign p2_smul_57596_comb = smul32b_32b_x_32b(p1_array_index_57048, p1_array_index_56956);
  assign p2_smul_57597_comb = smul32b_32b_x_32b(p1_array_index_57049, p1_array_index_56964);
  assign p2_smul_57598_comb = smul32b_32b_x_32b(p1_array_index_57050, p1_array_index_56962);
  assign p2_smul_57599_comb = smul32b_32b_x_32b(p1_array_index_57051, p1_array_index_56960);
  assign p2_smul_57600_comb = smul32b_32b_x_32b(p1_array_index_57052, p1_array_index_56958);
  assign p2_smul_57585_comb = smul32b_32b_x_32b(p1_array_index_57037, p1_array_index_57013);
  assign p2_smul_57586_comb = smul32b_32b_x_32b(p1_array_index_57038, p1_array_index_57014);
  assign p2_smul_57587_comb = smul32b_32b_x_32b(p1_array_index_57039, p1_array_index_57015);
  assign p2_smul_57588_comb = smul32b_32b_x_32b(p1_array_index_57040, p1_array_index_57016);
  assign p2_smul_57589_comb = smul32b_32b_x_32b(p1_array_index_57041, p1_array_index_57017);
  assign p2_smul_57590_comb = smul32b_32b_x_32b(p1_array_index_57042, p1_array_index_57018);
  assign p2_smul_57591_comb = smul32b_32b_x_32b(p1_array_index_57043, p1_array_index_57019);
  assign p2_smul_57592_comb = smul32b_32b_x_32b(p1_array_index_57044, p1_array_index_57020);
  assign p2_smul_57577_comb = smul32b_32b_x_32b(p1_array_index_57037, p1_array_index_57005);
  assign p2_smul_57578_comb = smul32b_32b_x_32b(p1_array_index_57038, p1_array_index_57006);
  assign p2_smul_57579_comb = smul32b_32b_x_32b(p1_array_index_57039, p1_array_index_57007);
  assign p2_smul_57580_comb = smul32b_32b_x_32b(p1_array_index_57040, p1_array_index_57008);
  assign p2_smul_57581_comb = smul32b_32b_x_32b(p1_array_index_57041, p1_array_index_57012);
  assign p2_smul_57582_comb = smul32b_32b_x_32b(p1_array_index_57042, p1_array_index_57011);
  assign p2_smul_57583_comb = smul32b_32b_x_32b(p1_array_index_57043, p1_array_index_57010);
  assign p2_smul_57584_comb = smul32b_32b_x_32b(p1_array_index_57044, p1_array_index_57009);
  assign p2_smul_57569_comb = smul32b_32b_x_32b(p1_array_index_57037, p1_array_index_56997);
  assign p2_smul_57570_comb = smul32b_32b_x_32b(p1_array_index_57038, p1_array_index_56998);
  assign p2_smul_57571_comb = smul32b_32b_x_32b(p1_array_index_57039, p1_array_index_56999);
  assign p2_smul_57572_comb = smul32b_32b_x_32b(p1_array_index_57040, p1_array_index_57000);
  assign p2_smul_57573_comb = smul32b_32b_x_32b(p1_array_index_57041, p1_array_index_57001);
  assign p2_smul_57574_comb = smul32b_32b_x_32b(p1_array_index_57042, p1_array_index_57002);
  assign p2_smul_57575_comb = smul32b_32b_x_32b(p1_array_index_57043, p1_array_index_57003);
  assign p2_smul_57576_comb = smul32b_32b_x_32b(p1_array_index_57044, p1_array_index_57004);
  assign p2_smul_57561_comb = smul32b_32b_x_32b(p1_array_index_57037, p1_array_index_56989);
  assign p2_smul_57562_comb = smul32b_32b_x_32b(p1_array_index_57038, p1_array_index_56990);
  assign p2_smul_57563_comb = smul32b_32b_x_32b(p1_array_index_57039, p1_array_index_56991);
  assign p2_smul_57564_comb = smul32b_32b_x_32b(p1_array_index_57040, p1_array_index_56992);
  assign p2_smul_57565_comb = smul32b_32b_x_32b(p1_array_index_57041, p1_array_index_56993);
  assign p2_smul_57566_comb = smul32b_32b_x_32b(p1_array_index_57042, p1_array_index_56994);
  assign p2_smul_57567_comb = smul32b_32b_x_32b(p1_array_index_57043, p1_array_index_56995);
  assign p2_smul_57568_comb = smul32b_32b_x_32b(p1_array_index_57044, p1_array_index_56996);
  assign p2_smul_57553_comb = smul32b_32b_x_32b(p1_array_index_57037, p1_array_index_56981);
  assign p2_smul_57554_comb = smul32b_32b_x_32b(p1_array_index_57038, p1_array_index_56982);
  assign p2_smul_57555_comb = smul32b_32b_x_32b(p1_array_index_57039, p1_array_index_56983);
  assign p2_smul_57556_comb = smul32b_32b_x_32b(p1_array_index_57040, p1_array_index_56984);
  assign p2_smul_57557_comb = smul32b_32b_x_32b(p1_array_index_57041, p1_array_index_56985);
  assign p2_smul_57558_comb = smul32b_32b_x_32b(p1_array_index_57042, p1_array_index_56986);
  assign p2_smul_57559_comb = smul32b_32b_x_32b(p1_array_index_57043, p1_array_index_56987);
  assign p2_smul_57560_comb = smul32b_32b_x_32b(p1_array_index_57044, p1_array_index_56988);
  assign p2_smul_57545_comb = smul32b_32b_x_32b(p1_array_index_57037, p1_array_index_56973);
  assign p2_smul_57546_comb = smul32b_32b_x_32b(p1_array_index_57038, p1_array_index_56974);
  assign p2_smul_57547_comb = smul32b_32b_x_32b(p1_array_index_57039, p1_array_index_56975);
  assign p2_smul_57548_comb = smul32b_32b_x_32b(p1_array_index_57040, p1_array_index_56976);
  assign p2_smul_57549_comb = smul32b_32b_x_32b(p1_array_index_57041, p1_array_index_56977);
  assign p2_smul_57550_comb = smul32b_32b_x_32b(p1_array_index_57042, p1_array_index_56978);
  assign p2_smul_57551_comb = smul32b_32b_x_32b(p1_array_index_57043, p1_array_index_56979);
  assign p2_smul_57552_comb = smul32b_32b_x_32b(p1_array_index_57044, p1_array_index_56980);
  assign p2_smul_57537_comb = smul32b_32b_x_32b(p1_array_index_57037, p1_array_index_56965);
  assign p2_smul_57538_comb = smul32b_32b_x_32b(p1_array_index_57038, p1_array_index_56966);
  assign p2_smul_57539_comb = smul32b_32b_x_32b(p1_array_index_57039, p1_array_index_56967);
  assign p2_smul_57540_comb = smul32b_32b_x_32b(p1_array_index_57040, p1_array_index_56968);
  assign p2_smul_57541_comb = smul32b_32b_x_32b(p1_array_index_57041, p1_array_index_56969);
  assign p2_smul_57542_comb = smul32b_32b_x_32b(p1_array_index_57042, p1_array_index_56970);
  assign p2_smul_57543_comb = smul32b_32b_x_32b(p1_array_index_57043, p1_array_index_56971);
  assign p2_smul_57544_comb = smul32b_32b_x_32b(p1_array_index_57044, p1_array_index_56972);
  assign p2_smul_57529_comb = smul32b_32b_x_32b(p1_array_index_57037, p1_array_index_56950);
  assign p2_smul_57530_comb = smul32b_32b_x_32b(p1_array_index_57038, p1_array_index_56952);
  assign p2_smul_57531_comb = smul32b_32b_x_32b(p1_array_index_57039, p1_array_index_56954);
  assign p2_smul_57532_comb = smul32b_32b_x_32b(p1_array_index_57040, p1_array_index_56956);
  assign p2_smul_57533_comb = smul32b_32b_x_32b(p1_array_index_57041, p1_array_index_56958);
  assign p2_smul_57534_comb = smul32b_32b_x_32b(p1_array_index_57042, p1_array_index_56960);
  assign p2_smul_57535_comb = smul32b_32b_x_32b(p1_array_index_57043, p1_array_index_56962);
  assign p2_smul_57536_comb = smul32b_32b_x_32b(p1_array_index_57044, p1_array_index_56964);
  assign p2_smul_57521_comb = smul32b_32b_x_32b(p1_array_index_57029, p1_array_index_57013);
  assign p2_smul_57522_comb = smul32b_32b_x_32b(p1_array_index_57030, p1_array_index_57014);
  assign p2_smul_57523_comb = smul32b_32b_x_32b(p1_array_index_57031, p1_array_index_57015);
  assign p2_smul_57524_comb = smul32b_32b_x_32b(p1_array_index_57032, p1_array_index_57016);
  assign p2_smul_57525_comb = smul32b_32b_x_32b(p1_array_index_57033, p1_array_index_57017);
  assign p2_smul_57526_comb = smul32b_32b_x_32b(p1_array_index_57034, p1_array_index_57018);
  assign p2_smul_57527_comb = smul32b_32b_x_32b(p1_array_index_57035, p1_array_index_57019);
  assign p2_smul_57528_comb = smul32b_32b_x_32b(p1_array_index_57036, p1_array_index_57020);
  assign p2_smul_57513_comb = smul32b_32b_x_32b(p1_array_index_57029, p1_array_index_57005);
  assign p2_smul_57514_comb = smul32b_32b_x_32b(p1_array_index_57030, p1_array_index_57006);
  assign p2_smul_57515_comb = smul32b_32b_x_32b(p1_array_index_57031, p1_array_index_57007);
  assign p2_smul_57516_comb = smul32b_32b_x_32b(p1_array_index_57032, p1_array_index_57008);
  assign p2_smul_57517_comb = smul32b_32b_x_32b(p1_array_index_57033, p1_array_index_57012);
  assign p2_smul_57518_comb = smul32b_32b_x_32b(p1_array_index_57034, p1_array_index_57011);
  assign p2_smul_57519_comb = smul32b_32b_x_32b(p1_array_index_57035, p1_array_index_57010);
  assign p2_smul_57520_comb = smul32b_32b_x_32b(p1_array_index_57036, p1_array_index_57009);
  assign p2_smul_57505_comb = smul32b_32b_x_32b(p1_array_index_57029, p1_array_index_56997);
  assign p2_smul_57506_comb = smul32b_32b_x_32b(p1_array_index_57030, p1_array_index_56998);
  assign p2_smul_57507_comb = smul32b_32b_x_32b(p1_array_index_57031, p1_array_index_56999);
  assign p2_smul_57508_comb = smul32b_32b_x_32b(p1_array_index_57032, p1_array_index_57000);
  assign p2_smul_57509_comb = smul32b_32b_x_32b(p1_array_index_57033, p1_array_index_57001);
  assign p2_smul_57510_comb = smul32b_32b_x_32b(p1_array_index_57034, p1_array_index_57002);
  assign p2_smul_57511_comb = smul32b_32b_x_32b(p1_array_index_57035, p1_array_index_57003);
  assign p2_smul_57512_comb = smul32b_32b_x_32b(p1_array_index_57036, p1_array_index_57004);
  assign p2_smul_57497_comb = smul32b_32b_x_32b(p1_array_index_57029, p1_array_index_56989);
  assign p2_smul_57498_comb = smul32b_32b_x_32b(p1_array_index_57030, p1_array_index_56990);
  assign p2_smul_57499_comb = smul32b_32b_x_32b(p1_array_index_57031, p1_array_index_56991);
  assign p2_smul_57500_comb = smul32b_32b_x_32b(p1_array_index_57032, p1_array_index_56992);
  assign p2_smul_57501_comb = smul32b_32b_x_32b(p1_array_index_57033, p1_array_index_56993);
  assign p2_smul_57502_comb = smul32b_32b_x_32b(p1_array_index_57034, p1_array_index_56994);
  assign p2_smul_57503_comb = smul32b_32b_x_32b(p1_array_index_57035, p1_array_index_56995);
  assign p2_smul_57504_comb = smul32b_32b_x_32b(p1_array_index_57036, p1_array_index_56996);
  assign p2_smul_57489_comb = smul32b_32b_x_32b(p1_array_index_57029, p1_array_index_56981);
  assign p2_smul_57490_comb = smul32b_32b_x_32b(p1_array_index_57030, p1_array_index_56982);
  assign p2_smul_57491_comb = smul32b_32b_x_32b(p1_array_index_57031, p1_array_index_56983);
  assign p2_smul_57492_comb = smul32b_32b_x_32b(p1_array_index_57032, p1_array_index_56984);
  assign p2_smul_57493_comb = smul32b_32b_x_32b(p1_array_index_57033, p1_array_index_56985);
  assign p2_smul_57494_comb = smul32b_32b_x_32b(p1_array_index_57034, p1_array_index_56986);
  assign p2_smul_57495_comb = smul32b_32b_x_32b(p1_array_index_57035, p1_array_index_56987);
  assign p2_smul_57496_comb = smul32b_32b_x_32b(p1_array_index_57036, p1_array_index_56988);
  assign p2_smul_57481_comb = smul32b_32b_x_32b(p1_array_index_57029, p1_array_index_56973);
  assign p2_smul_57482_comb = smul32b_32b_x_32b(p1_array_index_57030, p1_array_index_56974);
  assign p2_smul_57483_comb = smul32b_32b_x_32b(p1_array_index_57031, p1_array_index_56975);
  assign p2_smul_57484_comb = smul32b_32b_x_32b(p1_array_index_57032, p1_array_index_56976);
  assign p2_smul_57485_comb = smul32b_32b_x_32b(p1_array_index_57033, p1_array_index_56977);
  assign p2_smul_57486_comb = smul32b_32b_x_32b(p1_array_index_57034, p1_array_index_56978);
  assign p2_smul_57487_comb = smul32b_32b_x_32b(p1_array_index_57035, p1_array_index_56979);
  assign p2_smul_57488_comb = smul32b_32b_x_32b(p1_array_index_57036, p1_array_index_56980);
  assign p2_smul_57473_comb = smul32b_32b_x_32b(p1_array_index_57029, p1_array_index_56965);
  assign p2_smul_57474_comb = smul32b_32b_x_32b(p1_array_index_57030, p1_array_index_56966);
  assign p2_smul_57475_comb = smul32b_32b_x_32b(p1_array_index_57031, p1_array_index_56967);
  assign p2_smul_57476_comb = smul32b_32b_x_32b(p1_array_index_57032, p1_array_index_56968);
  assign p2_smul_57477_comb = smul32b_32b_x_32b(p1_array_index_57033, p1_array_index_56969);
  assign p2_smul_57478_comb = smul32b_32b_x_32b(p1_array_index_57034, p1_array_index_56970);
  assign p2_smul_57479_comb = smul32b_32b_x_32b(p1_array_index_57035, p1_array_index_56971);
  assign p2_smul_57480_comb = smul32b_32b_x_32b(p1_array_index_57036, p1_array_index_56972);
  assign p2_smul_57465_comb = smul32b_32b_x_32b(p1_array_index_57029, p1_array_index_56950);
  assign p2_smul_57466_comb = smul32b_32b_x_32b(p1_array_index_57030, p1_array_index_56952);
  assign p2_smul_57467_comb = smul32b_32b_x_32b(p1_array_index_57031, p1_array_index_56954);
  assign p2_smul_57468_comb = smul32b_32b_x_32b(p1_array_index_57032, p1_array_index_56956);
  assign p2_smul_57469_comb = smul32b_32b_x_32b(p1_array_index_57033, p1_array_index_56958);
  assign p2_smul_57470_comb = smul32b_32b_x_32b(p1_array_index_57034, p1_array_index_56960);
  assign p2_smul_57471_comb = smul32b_32b_x_32b(p1_array_index_57035, p1_array_index_56962);
  assign p2_smul_57472_comb = smul32b_32b_x_32b(p1_array_index_57036, p1_array_index_56964);
  assign p2_smul_57457_comb = smul32b_32b_x_32b(p1_array_index_57021, p1_array_index_57013);
  assign p2_smul_57458_comb = smul32b_32b_x_32b(p1_array_index_57022, p1_array_index_57014);
  assign p2_smul_57459_comb = smul32b_32b_x_32b(p1_array_index_57023, p1_array_index_57015);
  assign p2_smul_57460_comb = smul32b_32b_x_32b(p1_array_index_57024, p1_array_index_57016);
  assign p2_smul_57461_comb = smul32b_32b_x_32b(p1_array_index_57025, p1_array_index_57017);
  assign p2_smul_57462_comb = smul32b_32b_x_32b(p1_array_index_57026, p1_array_index_57018);
  assign p2_smul_57463_comb = smul32b_32b_x_32b(p1_array_index_57027, p1_array_index_57019);
  assign p2_smul_57464_comb = smul32b_32b_x_32b(p1_array_index_57028, p1_array_index_57020);
  assign p2_smul_57449_comb = smul32b_32b_x_32b(p1_array_index_57021, p1_array_index_57005);
  assign p2_smul_57450_comb = smul32b_32b_x_32b(p1_array_index_57022, p1_array_index_57006);
  assign p2_smul_57451_comb = smul32b_32b_x_32b(p1_array_index_57023, p1_array_index_57007);
  assign p2_smul_57452_comb = smul32b_32b_x_32b(p1_array_index_57024, p1_array_index_57008);
  assign p2_smul_57453_comb = smul32b_32b_x_32b(p1_array_index_57025, p1_array_index_57012);
  assign p2_smul_57454_comb = smul32b_32b_x_32b(p1_array_index_57026, p1_array_index_57011);
  assign p2_smul_57455_comb = smul32b_32b_x_32b(p1_array_index_57027, p1_array_index_57010);
  assign p2_smul_57456_comb = smul32b_32b_x_32b(p1_array_index_57028, p1_array_index_57009);
  assign p2_smul_57441_comb = smul32b_32b_x_32b(p1_array_index_57021, p1_array_index_56997);
  assign p2_smul_57442_comb = smul32b_32b_x_32b(p1_array_index_57022, p1_array_index_56998);
  assign p2_smul_57443_comb = smul32b_32b_x_32b(p1_array_index_57023, p1_array_index_56999);
  assign p2_smul_57444_comb = smul32b_32b_x_32b(p1_array_index_57024, p1_array_index_57000);
  assign p2_smul_57445_comb = smul32b_32b_x_32b(p1_array_index_57025, p1_array_index_57001);
  assign p2_smul_57446_comb = smul32b_32b_x_32b(p1_array_index_57026, p1_array_index_57002);
  assign p2_smul_57447_comb = smul32b_32b_x_32b(p1_array_index_57027, p1_array_index_57003);
  assign p2_smul_57448_comb = smul32b_32b_x_32b(p1_array_index_57028, p1_array_index_57004);
  assign p2_smul_57433_comb = smul32b_32b_x_32b(p1_array_index_57021, p1_array_index_56989);
  assign p2_smul_57434_comb = smul32b_32b_x_32b(p1_array_index_57022, p1_array_index_56990);
  assign p2_smul_57435_comb = smul32b_32b_x_32b(p1_array_index_57023, p1_array_index_56991);
  assign p2_smul_57436_comb = smul32b_32b_x_32b(p1_array_index_57024, p1_array_index_56992);
  assign p2_smul_57437_comb = smul32b_32b_x_32b(p1_array_index_57025, p1_array_index_56993);
  assign p2_smul_57438_comb = smul32b_32b_x_32b(p1_array_index_57026, p1_array_index_56994);
  assign p2_smul_57439_comb = smul32b_32b_x_32b(p1_array_index_57027, p1_array_index_56995);
  assign p2_smul_57440_comb = smul32b_32b_x_32b(p1_array_index_57028, p1_array_index_56996);
  assign p2_smul_57425_comb = smul32b_32b_x_32b(p1_array_index_57021, p1_array_index_56981);
  assign p2_smul_57426_comb = smul32b_32b_x_32b(p1_array_index_57022, p1_array_index_56982);
  assign p2_smul_57427_comb = smul32b_32b_x_32b(p1_array_index_57023, p1_array_index_56983);
  assign p2_smul_57428_comb = smul32b_32b_x_32b(p1_array_index_57024, p1_array_index_56984);
  assign p2_smul_57429_comb = smul32b_32b_x_32b(p1_array_index_57025, p1_array_index_56985);
  assign p2_smul_57430_comb = smul32b_32b_x_32b(p1_array_index_57026, p1_array_index_56986);
  assign p2_smul_57431_comb = smul32b_32b_x_32b(p1_array_index_57027, p1_array_index_56987);
  assign p2_smul_57432_comb = smul32b_32b_x_32b(p1_array_index_57028, p1_array_index_56988);
  assign p2_smul_57417_comb = smul32b_32b_x_32b(p1_array_index_57021, p1_array_index_56973);
  assign p2_smul_57418_comb = smul32b_32b_x_32b(p1_array_index_57022, p1_array_index_56974);
  assign p2_smul_57419_comb = smul32b_32b_x_32b(p1_array_index_57023, p1_array_index_56975);
  assign p2_smul_57420_comb = smul32b_32b_x_32b(p1_array_index_57024, p1_array_index_56976);
  assign p2_smul_57421_comb = smul32b_32b_x_32b(p1_array_index_57025, p1_array_index_56977);
  assign p2_smul_57422_comb = smul32b_32b_x_32b(p1_array_index_57026, p1_array_index_56978);
  assign p2_smul_57423_comb = smul32b_32b_x_32b(p1_array_index_57027, p1_array_index_56979);
  assign p2_smul_57424_comb = smul32b_32b_x_32b(p1_array_index_57028, p1_array_index_56980);
  assign p2_smul_57409_comb = smul32b_32b_x_32b(p1_array_index_57021, p1_array_index_56965);
  assign p2_smul_57410_comb = smul32b_32b_x_32b(p1_array_index_57022, p1_array_index_56966);
  assign p2_smul_57411_comb = smul32b_32b_x_32b(p1_array_index_57023, p1_array_index_56967);
  assign p2_smul_57412_comb = smul32b_32b_x_32b(p1_array_index_57024, p1_array_index_56968);
  assign p2_smul_57413_comb = smul32b_32b_x_32b(p1_array_index_57025, p1_array_index_56969);
  assign p2_smul_57414_comb = smul32b_32b_x_32b(p1_array_index_57026, p1_array_index_56970);
  assign p2_smul_57415_comb = smul32b_32b_x_32b(p1_array_index_57027, p1_array_index_56971);
  assign p2_smul_57416_comb = smul32b_32b_x_32b(p1_array_index_57028, p1_array_index_56972);
  assign p2_smul_57401_comb = smul32b_32b_x_32b(p1_array_index_57021, p1_array_index_56950);
  assign p2_smul_57402_comb = smul32b_32b_x_32b(p1_array_index_57022, p1_array_index_56952);
  assign p2_smul_57403_comb = smul32b_32b_x_32b(p1_array_index_57023, p1_array_index_56954);
  assign p2_smul_57404_comb = smul32b_32b_x_32b(p1_array_index_57024, p1_array_index_56956);
  assign p2_smul_57405_comb = smul32b_32b_x_32b(p1_array_index_57025, p1_array_index_56958);
  assign p2_smul_57406_comb = smul32b_32b_x_32b(p1_array_index_57026, p1_array_index_56960);
  assign p2_smul_57407_comb = smul32b_32b_x_32b(p1_array_index_57027, p1_array_index_56962);
  assign p2_smul_57408_comb = smul32b_32b_x_32b(p1_array_index_57028, p1_array_index_56964);
  assign p2_smul_57393_comb = smul32b_32b_x_32b(p1_array_index_56949, p1_array_index_57013);
  assign p2_smul_57394_comb = smul32b_32b_x_32b(p1_array_index_56951, p1_array_index_57014);
  assign p2_smul_57395_comb = smul32b_32b_x_32b(p1_array_index_56953, p1_array_index_57015);
  assign p2_smul_57396_comb = smul32b_32b_x_32b(p1_array_index_56955, p1_array_index_57016);
  assign p2_smul_57397_comb = smul32b_32b_x_32b(p1_array_index_56957, p1_array_index_57017);
  assign p2_smul_57398_comb = smul32b_32b_x_32b(p1_array_index_56959, p1_array_index_57018);
  assign p2_smul_57399_comb = smul32b_32b_x_32b(p1_array_index_56961, p1_array_index_57019);
  assign p2_smul_57400_comb = smul32b_32b_x_32b(p1_array_index_56963, p1_array_index_57020);
  assign p2_smul_57385_comb = smul32b_32b_x_32b(p1_array_index_56949, p1_array_index_57005);
  assign p2_smul_57386_comb = smul32b_32b_x_32b(p1_array_index_56951, p1_array_index_57006);
  assign p2_smul_57387_comb = smul32b_32b_x_32b(p1_array_index_56953, p1_array_index_57007);
  assign p2_smul_57388_comb = smul32b_32b_x_32b(p1_array_index_56955, p1_array_index_57008);
  assign p2_smul_57389_comb = smul32b_32b_x_32b(p1_array_index_56963, p1_array_index_57009);
  assign p2_smul_57390_comb = smul32b_32b_x_32b(p1_array_index_56961, p1_array_index_57010);
  assign p2_smul_57391_comb = smul32b_32b_x_32b(p1_array_index_56959, p1_array_index_57011);
  assign p2_smul_57392_comb = smul32b_32b_x_32b(p1_array_index_56957, p1_array_index_57012);
  assign p2_smul_57377_comb = smul32b_32b_x_32b(p1_array_index_56949, p1_array_index_56997);
  assign p2_smul_57378_comb = smul32b_32b_x_32b(p1_array_index_56951, p1_array_index_56998);
  assign p2_smul_57379_comb = smul32b_32b_x_32b(p1_array_index_56953, p1_array_index_56999);
  assign p2_smul_57380_comb = smul32b_32b_x_32b(p1_array_index_56955, p1_array_index_57000);
  assign p2_smul_57381_comb = smul32b_32b_x_32b(p1_array_index_56957, p1_array_index_57001);
  assign p2_smul_57382_comb = smul32b_32b_x_32b(p1_array_index_56959, p1_array_index_57002);
  assign p2_smul_57383_comb = smul32b_32b_x_32b(p1_array_index_56961, p1_array_index_57003);
  assign p2_smul_57384_comb = smul32b_32b_x_32b(p1_array_index_56963, p1_array_index_57004);
  assign p2_smul_57369_comb = smul32b_32b_x_32b(p1_array_index_56949, p1_array_index_56989);
  assign p2_smul_57370_comb = smul32b_32b_x_32b(p1_array_index_56951, p1_array_index_56990);
  assign p2_smul_57371_comb = smul32b_32b_x_32b(p1_array_index_56953, p1_array_index_56991);
  assign p2_smul_57372_comb = smul32b_32b_x_32b(p1_array_index_56955, p1_array_index_56992);
  assign p2_smul_57373_comb = smul32b_32b_x_32b(p1_array_index_56957, p1_array_index_56993);
  assign p2_smul_57374_comb = smul32b_32b_x_32b(p1_array_index_56959, p1_array_index_56994);
  assign p2_smul_57375_comb = smul32b_32b_x_32b(p1_array_index_56961, p1_array_index_56995);
  assign p2_smul_57376_comb = smul32b_32b_x_32b(p1_array_index_56963, p1_array_index_56996);
  assign p2_smul_57361_comb = smul32b_32b_x_32b(p1_array_index_56949, p1_array_index_56981);
  assign p2_smul_57362_comb = smul32b_32b_x_32b(p1_array_index_56951, p1_array_index_56982);
  assign p2_smul_57363_comb = smul32b_32b_x_32b(p1_array_index_56953, p1_array_index_56983);
  assign p2_smul_57364_comb = smul32b_32b_x_32b(p1_array_index_56955, p1_array_index_56984);
  assign p2_smul_57365_comb = smul32b_32b_x_32b(p1_array_index_56957, p1_array_index_56985);
  assign p2_smul_57366_comb = smul32b_32b_x_32b(p1_array_index_56959, p1_array_index_56986);
  assign p2_smul_57367_comb = smul32b_32b_x_32b(p1_array_index_56961, p1_array_index_56987);
  assign p2_smul_57368_comb = smul32b_32b_x_32b(p1_array_index_56963, p1_array_index_56988);
  assign p2_smul_57353_comb = smul32b_32b_x_32b(p1_array_index_56949, p1_array_index_56973);
  assign p2_smul_57354_comb = smul32b_32b_x_32b(p1_array_index_56951, p1_array_index_56974);
  assign p2_smul_57355_comb = smul32b_32b_x_32b(p1_array_index_56953, p1_array_index_56975);
  assign p2_smul_57356_comb = smul32b_32b_x_32b(p1_array_index_56955, p1_array_index_56976);
  assign p2_smul_57357_comb = smul32b_32b_x_32b(p1_array_index_56957, p1_array_index_56977);
  assign p2_smul_57358_comb = smul32b_32b_x_32b(p1_array_index_56959, p1_array_index_56978);
  assign p2_smul_57359_comb = smul32b_32b_x_32b(p1_array_index_56961, p1_array_index_56979);
  assign p2_smul_57360_comb = smul32b_32b_x_32b(p1_array_index_56963, p1_array_index_56980);
  assign p2_smul_57345_comb = smul32b_32b_x_32b(p1_array_index_56949, p1_array_index_56965);
  assign p2_smul_57346_comb = smul32b_32b_x_32b(p1_array_index_56951, p1_array_index_56966);
  assign p2_smul_57347_comb = smul32b_32b_x_32b(p1_array_index_56953, p1_array_index_56967);
  assign p2_smul_57348_comb = smul32b_32b_x_32b(p1_array_index_56955, p1_array_index_56968);
  assign p2_smul_57349_comb = smul32b_32b_x_32b(p1_array_index_56957, p1_array_index_56969);
  assign p2_smul_57350_comb = smul32b_32b_x_32b(p1_array_index_56959, p1_array_index_56970);
  assign p2_smul_57351_comb = smul32b_32b_x_32b(p1_array_index_56961, p1_array_index_56971);
  assign p2_smul_57352_comb = smul32b_32b_x_32b(p1_array_index_56963, p1_array_index_56972);
  assign p2_smul_57337_comb = smul32b_32b_x_32b(p1_array_index_56949, p1_array_index_56950);
  assign p2_smul_57338_comb = smul32b_32b_x_32b(p1_array_index_56951, p1_array_index_56952);
  assign p2_smul_57339_comb = smul32b_32b_x_32b(p1_array_index_56953, p1_array_index_56954);
  assign p2_smul_57340_comb = smul32b_32b_x_32b(p1_array_index_56955, p1_array_index_56956);
  assign p2_smul_57341_comb = smul32b_32b_x_32b(p1_array_index_56957, p1_array_index_56958);
  assign p2_smul_57342_comb = smul32b_32b_x_32b(p1_array_index_56959, p1_array_index_56960);
  assign p2_smul_57343_comb = smul32b_32b_x_32b(p1_array_index_56961, p1_array_index_56962);
  assign p2_smul_57344_comb = smul32b_32b_x_32b(p1_array_index_56963, p1_array_index_56964);
  assign p2_add_58101_comb = p2_smul_57841_comb + p2_smul_57842_comb;
  assign p2_add_58102_comb = p2_smul_57843_comb + p2_smul_57844_comb;
  assign p2_add_58103_comb = p2_smul_57845_comb + p2_smul_57846_comb;
  assign p2_add_58104_comb = p2_smul_57847_comb + p2_smul_57848_comb;
  assign p2_add_58097_comb = p2_smul_57833_comb + p2_smul_57834_comb;
  assign p2_add_58098_comb = p2_smul_57835_comb + p2_smul_57836_comb;
  assign p2_add_58099_comb = p2_smul_57837_comb + p2_smul_57838_comb;
  assign p2_add_58100_comb = p2_smul_57839_comb + p2_smul_57840_comb;
  assign p2_add_58093_comb = p2_smul_57825_comb + p2_smul_57826_comb;
  assign p2_add_58094_comb = p2_smul_57827_comb + p2_smul_57828_comb;
  assign p2_add_58095_comb = p2_smul_57829_comb + p2_smul_57830_comb;
  assign p2_add_58096_comb = p2_smul_57831_comb + p2_smul_57832_comb;
  assign p2_add_58089_comb = p2_smul_57817_comb + p2_smul_57818_comb;
  assign p2_add_58090_comb = p2_smul_57819_comb + p2_smul_57820_comb;
  assign p2_add_58091_comb = p2_smul_57821_comb + p2_smul_57822_comb;
  assign p2_add_58092_comb = p2_smul_57823_comb + p2_smul_57824_comb;
  assign p2_add_58085_comb = p2_smul_57809_comb + p2_smul_57810_comb;
  assign p2_add_58086_comb = p2_smul_57811_comb + p2_smul_57812_comb;
  assign p2_add_58087_comb = p2_smul_57813_comb + p2_smul_57814_comb;
  assign p2_add_58088_comb = p2_smul_57815_comb + p2_smul_57816_comb;
  assign p2_add_58081_comb = p2_smul_57801_comb + p2_smul_57802_comb;
  assign p2_add_58082_comb = p2_smul_57803_comb + p2_smul_57804_comb;
  assign p2_add_58083_comb = p2_smul_57805_comb + p2_smul_57806_comb;
  assign p2_add_58084_comb = p2_smul_57807_comb + p2_smul_57808_comb;
  assign p2_add_58077_comb = p2_smul_57793_comb + p2_smul_57794_comb;
  assign p2_add_58078_comb = p2_smul_57795_comb + p2_smul_57796_comb;
  assign p2_add_58079_comb = p2_smul_57797_comb + p2_smul_57798_comb;
  assign p2_add_58080_comb = p2_smul_57799_comb + p2_smul_57800_comb;
  assign p2_add_58073_comb = p2_smul_57785_comb + p2_smul_57786_comb;
  assign p2_add_58074_comb = p2_smul_57787_comb + p2_smul_57788_comb;
  assign p2_add_58075_comb = p2_smul_57789_comb + p2_smul_57790_comb;
  assign p2_add_58076_comb = p2_smul_57791_comb + p2_smul_57792_comb;
  assign p2_add_58069_comb = p2_smul_57777_comb + p2_smul_57778_comb;
  assign p2_add_58070_comb = p2_smul_57779_comb + p2_smul_57780_comb;
  assign p2_add_58071_comb = p2_smul_57781_comb + p2_smul_57782_comb;
  assign p2_add_58072_comb = p2_smul_57783_comb + p2_smul_57784_comb;
  assign p2_add_58065_comb = p2_smul_57769_comb + p2_smul_57770_comb;
  assign p2_add_58066_comb = p2_smul_57771_comb + p2_smul_57772_comb;
  assign p2_add_58067_comb = p2_smul_57773_comb + p2_smul_57774_comb;
  assign p2_add_58068_comb = p2_smul_57775_comb + p2_smul_57776_comb;
  assign p2_add_58061_comb = p2_smul_57761_comb + p2_smul_57762_comb;
  assign p2_add_58062_comb = p2_smul_57763_comb + p2_smul_57764_comb;
  assign p2_add_58063_comb = p2_smul_57765_comb + p2_smul_57766_comb;
  assign p2_add_58064_comb = p2_smul_57767_comb + p2_smul_57768_comb;
  assign p2_add_58057_comb = p2_smul_57753_comb + p2_smul_57754_comb;
  assign p2_add_58058_comb = p2_smul_57755_comb + p2_smul_57756_comb;
  assign p2_add_58059_comb = p2_smul_57757_comb + p2_smul_57758_comb;
  assign p2_add_58060_comb = p2_smul_57759_comb + p2_smul_57760_comb;
  assign p2_add_58053_comb = p2_smul_57745_comb + p2_smul_57746_comb;
  assign p2_add_58054_comb = p2_smul_57747_comb + p2_smul_57748_comb;
  assign p2_add_58055_comb = p2_smul_57749_comb + p2_smul_57750_comb;
  assign p2_add_58056_comb = p2_smul_57751_comb + p2_smul_57752_comb;
  assign p2_add_58049_comb = p2_smul_57737_comb + p2_smul_57738_comb;
  assign p2_add_58050_comb = p2_smul_57739_comb + p2_smul_57740_comb;
  assign p2_add_58051_comb = p2_smul_57741_comb + p2_smul_57742_comb;
  assign p2_add_58052_comb = p2_smul_57743_comb + p2_smul_57744_comb;
  assign p2_add_58045_comb = p2_smul_57729_comb + p2_smul_57730_comb;
  assign p2_add_58046_comb = p2_smul_57731_comb + p2_smul_57732_comb;
  assign p2_add_58047_comb = p2_smul_57733_comb + p2_smul_57734_comb;
  assign p2_add_58048_comb = p2_smul_57735_comb + p2_smul_57736_comb;
  assign p2_add_58041_comb = p2_smul_57721_comb + p2_smul_57722_comb;
  assign p2_add_58042_comb = p2_smul_57723_comb + p2_smul_57724_comb;
  assign p2_add_58043_comb = p2_smul_57725_comb + p2_smul_57726_comb;
  assign p2_add_58044_comb = p2_smul_57727_comb + p2_smul_57728_comb;
  assign p2_add_58037_comb = p2_smul_57713_comb + p2_smul_57714_comb;
  assign p2_add_58038_comb = p2_smul_57715_comb + p2_smul_57716_comb;
  assign p2_add_58039_comb = p2_smul_57717_comb + p2_smul_57718_comb;
  assign p2_add_58040_comb = p2_smul_57719_comb + p2_smul_57720_comb;
  assign p2_add_58033_comb = p2_smul_57705_comb + p2_smul_57706_comb;
  assign p2_add_58034_comb = p2_smul_57707_comb + p2_smul_57708_comb;
  assign p2_add_58035_comb = p2_smul_57709_comb + p2_smul_57710_comb;
  assign p2_add_58036_comb = p2_smul_57711_comb + p2_smul_57712_comb;
  assign p2_add_58029_comb = p2_smul_57697_comb + p2_smul_57698_comb;
  assign p2_add_58030_comb = p2_smul_57699_comb + p2_smul_57700_comb;
  assign p2_add_58031_comb = p2_smul_57701_comb + p2_smul_57702_comb;
  assign p2_add_58032_comb = p2_smul_57703_comb + p2_smul_57704_comb;
  assign p2_add_58025_comb = p2_smul_57689_comb + p2_smul_57690_comb;
  assign p2_add_58026_comb = p2_smul_57691_comb + p2_smul_57692_comb;
  assign p2_add_58027_comb = p2_smul_57693_comb + p2_smul_57694_comb;
  assign p2_add_58028_comb = p2_smul_57695_comb + p2_smul_57696_comb;
  assign p2_add_58021_comb = p2_smul_57681_comb + p2_smul_57682_comb;
  assign p2_add_58022_comb = p2_smul_57683_comb + p2_smul_57684_comb;
  assign p2_add_58023_comb = p2_smul_57685_comb + p2_smul_57686_comb;
  assign p2_add_58024_comb = p2_smul_57687_comb + p2_smul_57688_comb;
  assign p2_add_58017_comb = p2_smul_57673_comb + p2_smul_57674_comb;
  assign p2_add_58018_comb = p2_smul_57675_comb + p2_smul_57676_comb;
  assign p2_add_58019_comb = p2_smul_57677_comb + p2_smul_57678_comb;
  assign p2_add_58020_comb = p2_smul_57679_comb + p2_smul_57680_comb;
  assign p2_add_58013_comb = p2_smul_57665_comb + p2_smul_57666_comb;
  assign p2_add_58014_comb = p2_smul_57667_comb + p2_smul_57668_comb;
  assign p2_add_58015_comb = p2_smul_57669_comb + p2_smul_57670_comb;
  assign p2_add_58016_comb = p2_smul_57671_comb + p2_smul_57672_comb;
  assign p2_add_58009_comb = p2_smul_57657_comb + p2_smul_57658_comb;
  assign p2_add_58010_comb = p2_smul_57659_comb + p2_smul_57660_comb;
  assign p2_add_58011_comb = p2_smul_57661_comb + p2_smul_57662_comb;
  assign p2_add_58012_comb = p2_smul_57663_comb + p2_smul_57664_comb;
  assign p2_add_58005_comb = p2_smul_57649_comb + p2_smul_57650_comb;
  assign p2_add_58006_comb = p2_smul_57651_comb + p2_smul_57652_comb;
  assign p2_add_58007_comb = p2_smul_57653_comb + p2_smul_57654_comb;
  assign p2_add_58008_comb = p2_smul_57655_comb + p2_smul_57656_comb;
  assign p2_add_58001_comb = p2_smul_57641_comb + p2_smul_57642_comb;
  assign p2_add_58002_comb = p2_smul_57643_comb + p2_smul_57644_comb;
  assign p2_add_58003_comb = p2_smul_57645_comb + p2_smul_57646_comb;
  assign p2_add_58004_comb = p2_smul_57647_comb + p2_smul_57648_comb;
  assign p2_add_57997_comb = p2_smul_57633_comb + p2_smul_57634_comb;
  assign p2_add_57998_comb = p2_smul_57635_comb + p2_smul_57636_comb;
  assign p2_add_57999_comb = p2_smul_57637_comb + p2_smul_57638_comb;
  assign p2_add_58000_comb = p2_smul_57639_comb + p2_smul_57640_comb;
  assign p2_add_57993_comb = p2_smul_57625_comb + p2_smul_57626_comb;
  assign p2_add_57994_comb = p2_smul_57627_comb + p2_smul_57628_comb;
  assign p2_add_57995_comb = p2_smul_57629_comb + p2_smul_57630_comb;
  assign p2_add_57996_comb = p2_smul_57631_comb + p2_smul_57632_comb;
  assign p2_add_57989_comb = p2_smul_57617_comb + p2_smul_57618_comb;
  assign p2_add_57990_comb = p2_smul_57619_comb + p2_smul_57620_comb;
  assign p2_add_57991_comb = p2_smul_57621_comb + p2_smul_57622_comb;
  assign p2_add_57992_comb = p2_smul_57623_comb + p2_smul_57624_comb;
  assign p2_add_57985_comb = p2_smul_57609_comb + p2_smul_57610_comb;
  assign p2_add_57986_comb = p2_smul_57611_comb + p2_smul_57612_comb;
  assign p2_add_57987_comb = p2_smul_57613_comb + p2_smul_57614_comb;
  assign p2_add_57988_comb = p2_smul_57615_comb + p2_smul_57616_comb;
  assign p2_add_57981_comb = p2_smul_57601_comb + p2_smul_57602_comb;
  assign p2_add_57982_comb = p2_smul_57603_comb + p2_smul_57604_comb;
  assign p2_add_57983_comb = p2_smul_57605_comb + p2_smul_57606_comb;
  assign p2_add_57984_comb = p2_smul_57607_comb + p2_smul_57608_comb;
  assign p2_add_57977_comb = p2_smul_57593_comb + p2_smul_57594_comb;
  assign p2_add_57978_comb = p2_smul_57595_comb + p2_smul_57596_comb;
  assign p2_add_57979_comb = p2_smul_57597_comb + p2_smul_57598_comb;
  assign p2_add_57980_comb = p2_smul_57599_comb + p2_smul_57600_comb;
  assign p2_add_57973_comb = p2_smul_57585_comb + p2_smul_57586_comb;
  assign p2_add_57974_comb = p2_smul_57587_comb + p2_smul_57588_comb;
  assign p2_add_57975_comb = p2_smul_57589_comb + p2_smul_57590_comb;
  assign p2_add_57976_comb = p2_smul_57591_comb + p2_smul_57592_comb;
  assign p2_add_57969_comb = p2_smul_57577_comb + p2_smul_57578_comb;
  assign p2_add_57970_comb = p2_smul_57579_comb + p2_smul_57580_comb;
  assign p2_add_57971_comb = p2_smul_57581_comb + p2_smul_57582_comb;
  assign p2_add_57972_comb = p2_smul_57583_comb + p2_smul_57584_comb;
  assign p2_add_57965_comb = p2_smul_57569_comb + p2_smul_57570_comb;
  assign p2_add_57966_comb = p2_smul_57571_comb + p2_smul_57572_comb;
  assign p2_add_57967_comb = p2_smul_57573_comb + p2_smul_57574_comb;
  assign p2_add_57968_comb = p2_smul_57575_comb + p2_smul_57576_comb;
  assign p2_add_57961_comb = p2_smul_57561_comb + p2_smul_57562_comb;
  assign p2_add_57962_comb = p2_smul_57563_comb + p2_smul_57564_comb;
  assign p2_add_57963_comb = p2_smul_57565_comb + p2_smul_57566_comb;
  assign p2_add_57964_comb = p2_smul_57567_comb + p2_smul_57568_comb;
  assign p2_add_57957_comb = p2_smul_57553_comb + p2_smul_57554_comb;
  assign p2_add_57958_comb = p2_smul_57555_comb + p2_smul_57556_comb;
  assign p2_add_57959_comb = p2_smul_57557_comb + p2_smul_57558_comb;
  assign p2_add_57960_comb = p2_smul_57559_comb + p2_smul_57560_comb;
  assign p2_add_57953_comb = p2_smul_57545_comb + p2_smul_57546_comb;
  assign p2_add_57954_comb = p2_smul_57547_comb + p2_smul_57548_comb;
  assign p2_add_57955_comb = p2_smul_57549_comb + p2_smul_57550_comb;
  assign p2_add_57956_comb = p2_smul_57551_comb + p2_smul_57552_comb;
  assign p2_add_57949_comb = p2_smul_57537_comb + p2_smul_57538_comb;
  assign p2_add_57950_comb = p2_smul_57539_comb + p2_smul_57540_comb;
  assign p2_add_57951_comb = p2_smul_57541_comb + p2_smul_57542_comb;
  assign p2_add_57952_comb = p2_smul_57543_comb + p2_smul_57544_comb;
  assign p2_add_57945_comb = p2_smul_57529_comb + p2_smul_57530_comb;
  assign p2_add_57946_comb = p2_smul_57531_comb + p2_smul_57532_comb;
  assign p2_add_57947_comb = p2_smul_57533_comb + p2_smul_57534_comb;
  assign p2_add_57948_comb = p2_smul_57535_comb + p2_smul_57536_comb;
  assign p2_add_57941_comb = p2_smul_57521_comb + p2_smul_57522_comb;
  assign p2_add_57942_comb = p2_smul_57523_comb + p2_smul_57524_comb;
  assign p2_add_57943_comb = p2_smul_57525_comb + p2_smul_57526_comb;
  assign p2_add_57944_comb = p2_smul_57527_comb + p2_smul_57528_comb;
  assign p2_add_57937_comb = p2_smul_57513_comb + p2_smul_57514_comb;
  assign p2_add_57938_comb = p2_smul_57515_comb + p2_smul_57516_comb;
  assign p2_add_57939_comb = p2_smul_57517_comb + p2_smul_57518_comb;
  assign p2_add_57940_comb = p2_smul_57519_comb + p2_smul_57520_comb;
  assign p2_add_57933_comb = p2_smul_57505_comb + p2_smul_57506_comb;
  assign p2_add_57934_comb = p2_smul_57507_comb + p2_smul_57508_comb;
  assign p2_add_57935_comb = p2_smul_57509_comb + p2_smul_57510_comb;
  assign p2_add_57936_comb = p2_smul_57511_comb + p2_smul_57512_comb;
  assign p2_add_57929_comb = p2_smul_57497_comb + p2_smul_57498_comb;
  assign p2_add_57930_comb = p2_smul_57499_comb + p2_smul_57500_comb;
  assign p2_add_57931_comb = p2_smul_57501_comb + p2_smul_57502_comb;
  assign p2_add_57932_comb = p2_smul_57503_comb + p2_smul_57504_comb;
  assign p2_add_57925_comb = p2_smul_57489_comb + p2_smul_57490_comb;
  assign p2_add_57926_comb = p2_smul_57491_comb + p2_smul_57492_comb;
  assign p2_add_57927_comb = p2_smul_57493_comb + p2_smul_57494_comb;
  assign p2_add_57928_comb = p2_smul_57495_comb + p2_smul_57496_comb;
  assign p2_add_57921_comb = p2_smul_57481_comb + p2_smul_57482_comb;
  assign p2_add_57922_comb = p2_smul_57483_comb + p2_smul_57484_comb;
  assign p2_add_57923_comb = p2_smul_57485_comb + p2_smul_57486_comb;
  assign p2_add_57924_comb = p2_smul_57487_comb + p2_smul_57488_comb;
  assign p2_add_57917_comb = p2_smul_57473_comb + p2_smul_57474_comb;
  assign p2_add_57918_comb = p2_smul_57475_comb + p2_smul_57476_comb;
  assign p2_add_57919_comb = p2_smul_57477_comb + p2_smul_57478_comb;
  assign p2_add_57920_comb = p2_smul_57479_comb + p2_smul_57480_comb;
  assign p2_add_57913_comb = p2_smul_57465_comb + p2_smul_57466_comb;
  assign p2_add_57914_comb = p2_smul_57467_comb + p2_smul_57468_comb;
  assign p2_add_57915_comb = p2_smul_57469_comb + p2_smul_57470_comb;
  assign p2_add_57916_comb = p2_smul_57471_comb + p2_smul_57472_comb;
  assign p2_add_57909_comb = p2_smul_57457_comb + p2_smul_57458_comb;
  assign p2_add_57910_comb = p2_smul_57459_comb + p2_smul_57460_comb;
  assign p2_add_57911_comb = p2_smul_57461_comb + p2_smul_57462_comb;
  assign p2_add_57912_comb = p2_smul_57463_comb + p2_smul_57464_comb;
  assign p2_add_57905_comb = p2_smul_57449_comb + p2_smul_57450_comb;
  assign p2_add_57906_comb = p2_smul_57451_comb + p2_smul_57452_comb;
  assign p2_add_57907_comb = p2_smul_57453_comb + p2_smul_57454_comb;
  assign p2_add_57908_comb = p2_smul_57455_comb + p2_smul_57456_comb;
  assign p2_add_57901_comb = p2_smul_57441_comb + p2_smul_57442_comb;
  assign p2_add_57902_comb = p2_smul_57443_comb + p2_smul_57444_comb;
  assign p2_add_57903_comb = p2_smul_57445_comb + p2_smul_57446_comb;
  assign p2_add_57904_comb = p2_smul_57447_comb + p2_smul_57448_comb;
  assign p2_add_57897_comb = p2_smul_57433_comb + p2_smul_57434_comb;
  assign p2_add_57898_comb = p2_smul_57435_comb + p2_smul_57436_comb;
  assign p2_add_57899_comb = p2_smul_57437_comb + p2_smul_57438_comb;
  assign p2_add_57900_comb = p2_smul_57439_comb + p2_smul_57440_comb;
  assign p2_add_57893_comb = p2_smul_57425_comb + p2_smul_57426_comb;
  assign p2_add_57894_comb = p2_smul_57427_comb + p2_smul_57428_comb;
  assign p2_add_57895_comb = p2_smul_57429_comb + p2_smul_57430_comb;
  assign p2_add_57896_comb = p2_smul_57431_comb + p2_smul_57432_comb;
  assign p2_add_57889_comb = p2_smul_57417_comb + p2_smul_57418_comb;
  assign p2_add_57890_comb = p2_smul_57419_comb + p2_smul_57420_comb;
  assign p2_add_57891_comb = p2_smul_57421_comb + p2_smul_57422_comb;
  assign p2_add_57892_comb = p2_smul_57423_comb + p2_smul_57424_comb;
  assign p2_add_57885_comb = p2_smul_57409_comb + p2_smul_57410_comb;
  assign p2_add_57886_comb = p2_smul_57411_comb + p2_smul_57412_comb;
  assign p2_add_57887_comb = p2_smul_57413_comb + p2_smul_57414_comb;
  assign p2_add_57888_comb = p2_smul_57415_comb + p2_smul_57416_comb;
  assign p2_add_57881_comb = p2_smul_57401_comb + p2_smul_57402_comb;
  assign p2_add_57882_comb = p2_smul_57403_comb + p2_smul_57404_comb;
  assign p2_add_57883_comb = p2_smul_57405_comb + p2_smul_57406_comb;
  assign p2_add_57884_comb = p2_smul_57407_comb + p2_smul_57408_comb;
  assign p2_add_57877_comb = p2_smul_57393_comb + p2_smul_57394_comb;
  assign p2_add_57878_comb = p2_smul_57395_comb + p2_smul_57396_comb;
  assign p2_add_57879_comb = p2_smul_57397_comb + p2_smul_57398_comb;
  assign p2_add_57880_comb = p2_smul_57399_comb + p2_smul_57400_comb;
  assign p2_add_57873_comb = p2_smul_57385_comb + p2_smul_57386_comb;
  assign p2_add_57874_comb = p2_smul_57387_comb + p2_smul_57388_comb;
  assign p2_add_57875_comb = p2_smul_57389_comb + p2_smul_57390_comb;
  assign p2_add_57876_comb = p2_smul_57391_comb + p2_smul_57392_comb;
  assign p2_add_57869_comb = p2_smul_57377_comb + p2_smul_57378_comb;
  assign p2_add_57870_comb = p2_smul_57379_comb + p2_smul_57380_comb;
  assign p2_add_57871_comb = p2_smul_57381_comb + p2_smul_57382_comb;
  assign p2_add_57872_comb = p2_smul_57383_comb + p2_smul_57384_comb;
  assign p2_add_57865_comb = p2_smul_57369_comb + p2_smul_57370_comb;
  assign p2_add_57866_comb = p2_smul_57371_comb + p2_smul_57372_comb;
  assign p2_add_57867_comb = p2_smul_57373_comb + p2_smul_57374_comb;
  assign p2_add_57868_comb = p2_smul_57375_comb + p2_smul_57376_comb;
  assign p2_add_57861_comb = p2_smul_57361_comb + p2_smul_57362_comb;
  assign p2_add_57862_comb = p2_smul_57363_comb + p2_smul_57364_comb;
  assign p2_add_57863_comb = p2_smul_57365_comb + p2_smul_57366_comb;
  assign p2_add_57864_comb = p2_smul_57367_comb + p2_smul_57368_comb;
  assign p2_add_57857_comb = p2_smul_57353_comb + p2_smul_57354_comb;
  assign p2_add_57858_comb = p2_smul_57355_comb + p2_smul_57356_comb;
  assign p2_add_57859_comb = p2_smul_57357_comb + p2_smul_57358_comb;
  assign p2_add_57860_comb = p2_smul_57359_comb + p2_smul_57360_comb;
  assign p2_add_57853_comb = p2_smul_57345_comb + p2_smul_57346_comb;
  assign p2_add_57854_comb = p2_smul_57347_comb + p2_smul_57348_comb;
  assign p2_add_57855_comb = p2_smul_57349_comb + p2_smul_57350_comb;
  assign p2_add_57856_comb = p2_smul_57351_comb + p2_smul_57352_comb;
  assign p2_add_57849_comb = p2_smul_57337_comb + p2_smul_57338_comb;
  assign p2_add_57850_comb = p2_smul_57339_comb + p2_smul_57340_comb;
  assign p2_add_57851_comb = p2_smul_57341_comb + p2_smul_57342_comb;
  assign p2_add_57852_comb = p2_smul_57343_comb + p2_smul_57344_comb;

  // Registers for pipe stage 2:
  reg [31:0] p2_a[8][8];
  reg [31:0] p2_b[8][8];
  reg [31:0] p2_add_58101;
  reg [31:0] p2_add_58102;
  reg [31:0] p2_add_58103;
  reg [31:0] p2_add_58104;
  reg [31:0] p2_add_58097;
  reg [31:0] p2_add_58098;
  reg [31:0] p2_add_58099;
  reg [31:0] p2_add_58100;
  reg [31:0] p2_add_58093;
  reg [31:0] p2_add_58094;
  reg [31:0] p2_add_58095;
  reg [31:0] p2_add_58096;
  reg [31:0] p2_add_58089;
  reg [31:0] p2_add_58090;
  reg [31:0] p2_add_58091;
  reg [31:0] p2_add_58092;
  reg [31:0] p2_add_58085;
  reg [31:0] p2_add_58086;
  reg [31:0] p2_add_58087;
  reg [31:0] p2_add_58088;
  reg [31:0] p2_add_58081;
  reg [31:0] p2_add_58082;
  reg [31:0] p2_add_58083;
  reg [31:0] p2_add_58084;
  reg [31:0] p2_add_58077;
  reg [31:0] p2_add_58078;
  reg [31:0] p2_add_58079;
  reg [31:0] p2_add_58080;
  reg [31:0] p2_add_58073;
  reg [31:0] p2_add_58074;
  reg [31:0] p2_add_58075;
  reg [31:0] p2_add_58076;
  reg [31:0] p2_add_58069;
  reg [31:0] p2_add_58070;
  reg [31:0] p2_add_58071;
  reg [31:0] p2_add_58072;
  reg [31:0] p2_add_58065;
  reg [31:0] p2_add_58066;
  reg [31:0] p2_add_58067;
  reg [31:0] p2_add_58068;
  reg [31:0] p2_add_58061;
  reg [31:0] p2_add_58062;
  reg [31:0] p2_add_58063;
  reg [31:0] p2_add_58064;
  reg [31:0] p2_add_58057;
  reg [31:0] p2_add_58058;
  reg [31:0] p2_add_58059;
  reg [31:0] p2_add_58060;
  reg [31:0] p2_add_58053;
  reg [31:0] p2_add_58054;
  reg [31:0] p2_add_58055;
  reg [31:0] p2_add_58056;
  reg [31:0] p2_add_58049;
  reg [31:0] p2_add_58050;
  reg [31:0] p2_add_58051;
  reg [31:0] p2_add_58052;
  reg [31:0] p2_add_58045;
  reg [31:0] p2_add_58046;
  reg [31:0] p2_add_58047;
  reg [31:0] p2_add_58048;
  reg [31:0] p2_add_58041;
  reg [31:0] p2_add_58042;
  reg [31:0] p2_add_58043;
  reg [31:0] p2_add_58044;
  reg [31:0] p2_add_58037;
  reg [31:0] p2_add_58038;
  reg [31:0] p2_add_58039;
  reg [31:0] p2_add_58040;
  reg [31:0] p2_add_58033;
  reg [31:0] p2_add_58034;
  reg [31:0] p2_add_58035;
  reg [31:0] p2_add_58036;
  reg [31:0] p2_add_58029;
  reg [31:0] p2_add_58030;
  reg [31:0] p2_add_58031;
  reg [31:0] p2_add_58032;
  reg [31:0] p2_add_58025;
  reg [31:0] p2_add_58026;
  reg [31:0] p2_add_58027;
  reg [31:0] p2_add_58028;
  reg [31:0] p2_add_58021;
  reg [31:0] p2_add_58022;
  reg [31:0] p2_add_58023;
  reg [31:0] p2_add_58024;
  reg [31:0] p2_add_58017;
  reg [31:0] p2_add_58018;
  reg [31:0] p2_add_58019;
  reg [31:0] p2_add_58020;
  reg [31:0] p2_add_58013;
  reg [31:0] p2_add_58014;
  reg [31:0] p2_add_58015;
  reg [31:0] p2_add_58016;
  reg [31:0] p2_add_58009;
  reg [31:0] p2_add_58010;
  reg [31:0] p2_add_58011;
  reg [31:0] p2_add_58012;
  reg [31:0] p2_add_58005;
  reg [31:0] p2_add_58006;
  reg [31:0] p2_add_58007;
  reg [31:0] p2_add_58008;
  reg [31:0] p2_add_58001;
  reg [31:0] p2_add_58002;
  reg [31:0] p2_add_58003;
  reg [31:0] p2_add_58004;
  reg [31:0] p2_add_57997;
  reg [31:0] p2_add_57998;
  reg [31:0] p2_add_57999;
  reg [31:0] p2_add_58000;
  reg [31:0] p2_add_57993;
  reg [31:0] p2_add_57994;
  reg [31:0] p2_add_57995;
  reg [31:0] p2_add_57996;
  reg [31:0] p2_add_57989;
  reg [31:0] p2_add_57990;
  reg [31:0] p2_add_57991;
  reg [31:0] p2_add_57992;
  reg [31:0] p2_add_57985;
  reg [31:0] p2_add_57986;
  reg [31:0] p2_add_57987;
  reg [31:0] p2_add_57988;
  reg [31:0] p2_add_57981;
  reg [31:0] p2_add_57982;
  reg [31:0] p2_add_57983;
  reg [31:0] p2_add_57984;
  reg [31:0] p2_add_57977;
  reg [31:0] p2_add_57978;
  reg [31:0] p2_add_57979;
  reg [31:0] p2_add_57980;
  reg [31:0] p2_add_57973;
  reg [31:0] p2_add_57974;
  reg [31:0] p2_add_57975;
  reg [31:0] p2_add_57976;
  reg [31:0] p2_add_57969;
  reg [31:0] p2_add_57970;
  reg [31:0] p2_add_57971;
  reg [31:0] p2_add_57972;
  reg [31:0] p2_add_57965;
  reg [31:0] p2_add_57966;
  reg [31:0] p2_add_57967;
  reg [31:0] p2_add_57968;
  reg [31:0] p2_add_57961;
  reg [31:0] p2_add_57962;
  reg [31:0] p2_add_57963;
  reg [31:0] p2_add_57964;
  reg [31:0] p2_add_57957;
  reg [31:0] p2_add_57958;
  reg [31:0] p2_add_57959;
  reg [31:0] p2_add_57960;
  reg [31:0] p2_add_57953;
  reg [31:0] p2_add_57954;
  reg [31:0] p2_add_57955;
  reg [31:0] p2_add_57956;
  reg [31:0] p2_add_57949;
  reg [31:0] p2_add_57950;
  reg [31:0] p2_add_57951;
  reg [31:0] p2_add_57952;
  reg [31:0] p2_add_57945;
  reg [31:0] p2_add_57946;
  reg [31:0] p2_add_57947;
  reg [31:0] p2_add_57948;
  reg [31:0] p2_add_57941;
  reg [31:0] p2_add_57942;
  reg [31:0] p2_add_57943;
  reg [31:0] p2_add_57944;
  reg [31:0] p2_add_57937;
  reg [31:0] p2_add_57938;
  reg [31:0] p2_add_57939;
  reg [31:0] p2_add_57940;
  reg [31:0] p2_add_57933;
  reg [31:0] p2_add_57934;
  reg [31:0] p2_add_57935;
  reg [31:0] p2_add_57936;
  reg [31:0] p2_add_57929;
  reg [31:0] p2_add_57930;
  reg [31:0] p2_add_57931;
  reg [31:0] p2_add_57932;
  reg [31:0] p2_add_57925;
  reg [31:0] p2_add_57926;
  reg [31:0] p2_add_57927;
  reg [31:0] p2_add_57928;
  reg [31:0] p2_add_57921;
  reg [31:0] p2_add_57922;
  reg [31:0] p2_add_57923;
  reg [31:0] p2_add_57924;
  reg [31:0] p2_add_57917;
  reg [31:0] p2_add_57918;
  reg [31:0] p2_add_57919;
  reg [31:0] p2_add_57920;
  reg [31:0] p2_add_57913;
  reg [31:0] p2_add_57914;
  reg [31:0] p2_add_57915;
  reg [31:0] p2_add_57916;
  reg [31:0] p2_add_57909;
  reg [31:0] p2_add_57910;
  reg [31:0] p2_add_57911;
  reg [31:0] p2_add_57912;
  reg [31:0] p2_add_57905;
  reg [31:0] p2_add_57906;
  reg [31:0] p2_add_57907;
  reg [31:0] p2_add_57908;
  reg [31:0] p2_add_57901;
  reg [31:0] p2_add_57902;
  reg [31:0] p2_add_57903;
  reg [31:0] p2_add_57904;
  reg [31:0] p2_add_57897;
  reg [31:0] p2_add_57898;
  reg [31:0] p2_add_57899;
  reg [31:0] p2_add_57900;
  reg [31:0] p2_add_57893;
  reg [31:0] p2_add_57894;
  reg [31:0] p2_add_57895;
  reg [31:0] p2_add_57896;
  reg [31:0] p2_add_57889;
  reg [31:0] p2_add_57890;
  reg [31:0] p2_add_57891;
  reg [31:0] p2_add_57892;
  reg [31:0] p2_add_57885;
  reg [31:0] p2_add_57886;
  reg [31:0] p2_add_57887;
  reg [31:0] p2_add_57888;
  reg [31:0] p2_add_57881;
  reg [31:0] p2_add_57882;
  reg [31:0] p2_add_57883;
  reg [31:0] p2_add_57884;
  reg [31:0] p2_add_57877;
  reg [31:0] p2_add_57878;
  reg [31:0] p2_add_57879;
  reg [31:0] p2_add_57880;
  reg [31:0] p2_add_57873;
  reg [31:0] p2_add_57874;
  reg [31:0] p2_add_57875;
  reg [31:0] p2_add_57876;
  reg [31:0] p2_add_57869;
  reg [31:0] p2_add_57870;
  reg [31:0] p2_add_57871;
  reg [31:0] p2_add_57872;
  reg [31:0] p2_add_57865;
  reg [31:0] p2_add_57866;
  reg [31:0] p2_add_57867;
  reg [31:0] p2_add_57868;
  reg [31:0] p2_add_57861;
  reg [31:0] p2_add_57862;
  reg [31:0] p2_add_57863;
  reg [31:0] p2_add_57864;
  reg [31:0] p2_add_57857;
  reg [31:0] p2_add_57858;
  reg [31:0] p2_add_57859;
  reg [31:0] p2_add_57860;
  reg [31:0] p2_add_57853;
  reg [31:0] p2_add_57854;
  reg [31:0] p2_add_57855;
  reg [31:0] p2_add_57856;
  reg [31:0] p2_add_57849;
  reg [31:0] p2_add_57850;
  reg [31:0] p2_add_57851;
  reg [31:0] p2_add_57852;
  always_ff @ (posedge clk) begin
    p2_a <= p1_a;
    p2_b <= p1_b;
    p2_add_58101 <= p2_add_58101_comb;
    p2_add_58102 <= p2_add_58102_comb;
    p2_add_58103 <= p2_add_58103_comb;
    p2_add_58104 <= p2_add_58104_comb;
    p2_add_58097 <= p2_add_58097_comb;
    p2_add_58098 <= p2_add_58098_comb;
    p2_add_58099 <= p2_add_58099_comb;
    p2_add_58100 <= p2_add_58100_comb;
    p2_add_58093 <= p2_add_58093_comb;
    p2_add_58094 <= p2_add_58094_comb;
    p2_add_58095 <= p2_add_58095_comb;
    p2_add_58096 <= p2_add_58096_comb;
    p2_add_58089 <= p2_add_58089_comb;
    p2_add_58090 <= p2_add_58090_comb;
    p2_add_58091 <= p2_add_58091_comb;
    p2_add_58092 <= p2_add_58092_comb;
    p2_add_58085 <= p2_add_58085_comb;
    p2_add_58086 <= p2_add_58086_comb;
    p2_add_58087 <= p2_add_58087_comb;
    p2_add_58088 <= p2_add_58088_comb;
    p2_add_58081 <= p2_add_58081_comb;
    p2_add_58082 <= p2_add_58082_comb;
    p2_add_58083 <= p2_add_58083_comb;
    p2_add_58084 <= p2_add_58084_comb;
    p2_add_58077 <= p2_add_58077_comb;
    p2_add_58078 <= p2_add_58078_comb;
    p2_add_58079 <= p2_add_58079_comb;
    p2_add_58080 <= p2_add_58080_comb;
    p2_add_58073 <= p2_add_58073_comb;
    p2_add_58074 <= p2_add_58074_comb;
    p2_add_58075 <= p2_add_58075_comb;
    p2_add_58076 <= p2_add_58076_comb;
    p2_add_58069 <= p2_add_58069_comb;
    p2_add_58070 <= p2_add_58070_comb;
    p2_add_58071 <= p2_add_58071_comb;
    p2_add_58072 <= p2_add_58072_comb;
    p2_add_58065 <= p2_add_58065_comb;
    p2_add_58066 <= p2_add_58066_comb;
    p2_add_58067 <= p2_add_58067_comb;
    p2_add_58068 <= p2_add_58068_comb;
    p2_add_58061 <= p2_add_58061_comb;
    p2_add_58062 <= p2_add_58062_comb;
    p2_add_58063 <= p2_add_58063_comb;
    p2_add_58064 <= p2_add_58064_comb;
    p2_add_58057 <= p2_add_58057_comb;
    p2_add_58058 <= p2_add_58058_comb;
    p2_add_58059 <= p2_add_58059_comb;
    p2_add_58060 <= p2_add_58060_comb;
    p2_add_58053 <= p2_add_58053_comb;
    p2_add_58054 <= p2_add_58054_comb;
    p2_add_58055 <= p2_add_58055_comb;
    p2_add_58056 <= p2_add_58056_comb;
    p2_add_58049 <= p2_add_58049_comb;
    p2_add_58050 <= p2_add_58050_comb;
    p2_add_58051 <= p2_add_58051_comb;
    p2_add_58052 <= p2_add_58052_comb;
    p2_add_58045 <= p2_add_58045_comb;
    p2_add_58046 <= p2_add_58046_comb;
    p2_add_58047 <= p2_add_58047_comb;
    p2_add_58048 <= p2_add_58048_comb;
    p2_add_58041 <= p2_add_58041_comb;
    p2_add_58042 <= p2_add_58042_comb;
    p2_add_58043 <= p2_add_58043_comb;
    p2_add_58044 <= p2_add_58044_comb;
    p2_add_58037 <= p2_add_58037_comb;
    p2_add_58038 <= p2_add_58038_comb;
    p2_add_58039 <= p2_add_58039_comb;
    p2_add_58040 <= p2_add_58040_comb;
    p2_add_58033 <= p2_add_58033_comb;
    p2_add_58034 <= p2_add_58034_comb;
    p2_add_58035 <= p2_add_58035_comb;
    p2_add_58036 <= p2_add_58036_comb;
    p2_add_58029 <= p2_add_58029_comb;
    p2_add_58030 <= p2_add_58030_comb;
    p2_add_58031 <= p2_add_58031_comb;
    p2_add_58032 <= p2_add_58032_comb;
    p2_add_58025 <= p2_add_58025_comb;
    p2_add_58026 <= p2_add_58026_comb;
    p2_add_58027 <= p2_add_58027_comb;
    p2_add_58028 <= p2_add_58028_comb;
    p2_add_58021 <= p2_add_58021_comb;
    p2_add_58022 <= p2_add_58022_comb;
    p2_add_58023 <= p2_add_58023_comb;
    p2_add_58024 <= p2_add_58024_comb;
    p2_add_58017 <= p2_add_58017_comb;
    p2_add_58018 <= p2_add_58018_comb;
    p2_add_58019 <= p2_add_58019_comb;
    p2_add_58020 <= p2_add_58020_comb;
    p2_add_58013 <= p2_add_58013_comb;
    p2_add_58014 <= p2_add_58014_comb;
    p2_add_58015 <= p2_add_58015_comb;
    p2_add_58016 <= p2_add_58016_comb;
    p2_add_58009 <= p2_add_58009_comb;
    p2_add_58010 <= p2_add_58010_comb;
    p2_add_58011 <= p2_add_58011_comb;
    p2_add_58012 <= p2_add_58012_comb;
    p2_add_58005 <= p2_add_58005_comb;
    p2_add_58006 <= p2_add_58006_comb;
    p2_add_58007 <= p2_add_58007_comb;
    p2_add_58008 <= p2_add_58008_comb;
    p2_add_58001 <= p2_add_58001_comb;
    p2_add_58002 <= p2_add_58002_comb;
    p2_add_58003 <= p2_add_58003_comb;
    p2_add_58004 <= p2_add_58004_comb;
    p2_add_57997 <= p2_add_57997_comb;
    p2_add_57998 <= p2_add_57998_comb;
    p2_add_57999 <= p2_add_57999_comb;
    p2_add_58000 <= p2_add_58000_comb;
    p2_add_57993 <= p2_add_57993_comb;
    p2_add_57994 <= p2_add_57994_comb;
    p2_add_57995 <= p2_add_57995_comb;
    p2_add_57996 <= p2_add_57996_comb;
    p2_add_57989 <= p2_add_57989_comb;
    p2_add_57990 <= p2_add_57990_comb;
    p2_add_57991 <= p2_add_57991_comb;
    p2_add_57992 <= p2_add_57992_comb;
    p2_add_57985 <= p2_add_57985_comb;
    p2_add_57986 <= p2_add_57986_comb;
    p2_add_57987 <= p2_add_57987_comb;
    p2_add_57988 <= p2_add_57988_comb;
    p2_add_57981 <= p2_add_57981_comb;
    p2_add_57982 <= p2_add_57982_comb;
    p2_add_57983 <= p2_add_57983_comb;
    p2_add_57984 <= p2_add_57984_comb;
    p2_add_57977 <= p2_add_57977_comb;
    p2_add_57978 <= p2_add_57978_comb;
    p2_add_57979 <= p2_add_57979_comb;
    p2_add_57980 <= p2_add_57980_comb;
    p2_add_57973 <= p2_add_57973_comb;
    p2_add_57974 <= p2_add_57974_comb;
    p2_add_57975 <= p2_add_57975_comb;
    p2_add_57976 <= p2_add_57976_comb;
    p2_add_57969 <= p2_add_57969_comb;
    p2_add_57970 <= p2_add_57970_comb;
    p2_add_57971 <= p2_add_57971_comb;
    p2_add_57972 <= p2_add_57972_comb;
    p2_add_57965 <= p2_add_57965_comb;
    p2_add_57966 <= p2_add_57966_comb;
    p2_add_57967 <= p2_add_57967_comb;
    p2_add_57968 <= p2_add_57968_comb;
    p2_add_57961 <= p2_add_57961_comb;
    p2_add_57962 <= p2_add_57962_comb;
    p2_add_57963 <= p2_add_57963_comb;
    p2_add_57964 <= p2_add_57964_comb;
    p2_add_57957 <= p2_add_57957_comb;
    p2_add_57958 <= p2_add_57958_comb;
    p2_add_57959 <= p2_add_57959_comb;
    p2_add_57960 <= p2_add_57960_comb;
    p2_add_57953 <= p2_add_57953_comb;
    p2_add_57954 <= p2_add_57954_comb;
    p2_add_57955 <= p2_add_57955_comb;
    p2_add_57956 <= p2_add_57956_comb;
    p2_add_57949 <= p2_add_57949_comb;
    p2_add_57950 <= p2_add_57950_comb;
    p2_add_57951 <= p2_add_57951_comb;
    p2_add_57952 <= p2_add_57952_comb;
    p2_add_57945 <= p2_add_57945_comb;
    p2_add_57946 <= p2_add_57946_comb;
    p2_add_57947 <= p2_add_57947_comb;
    p2_add_57948 <= p2_add_57948_comb;
    p2_add_57941 <= p2_add_57941_comb;
    p2_add_57942 <= p2_add_57942_comb;
    p2_add_57943 <= p2_add_57943_comb;
    p2_add_57944 <= p2_add_57944_comb;
    p2_add_57937 <= p2_add_57937_comb;
    p2_add_57938 <= p2_add_57938_comb;
    p2_add_57939 <= p2_add_57939_comb;
    p2_add_57940 <= p2_add_57940_comb;
    p2_add_57933 <= p2_add_57933_comb;
    p2_add_57934 <= p2_add_57934_comb;
    p2_add_57935 <= p2_add_57935_comb;
    p2_add_57936 <= p2_add_57936_comb;
    p2_add_57929 <= p2_add_57929_comb;
    p2_add_57930 <= p2_add_57930_comb;
    p2_add_57931 <= p2_add_57931_comb;
    p2_add_57932 <= p2_add_57932_comb;
    p2_add_57925 <= p2_add_57925_comb;
    p2_add_57926 <= p2_add_57926_comb;
    p2_add_57927 <= p2_add_57927_comb;
    p2_add_57928 <= p2_add_57928_comb;
    p2_add_57921 <= p2_add_57921_comb;
    p2_add_57922 <= p2_add_57922_comb;
    p2_add_57923 <= p2_add_57923_comb;
    p2_add_57924 <= p2_add_57924_comb;
    p2_add_57917 <= p2_add_57917_comb;
    p2_add_57918 <= p2_add_57918_comb;
    p2_add_57919 <= p2_add_57919_comb;
    p2_add_57920 <= p2_add_57920_comb;
    p2_add_57913 <= p2_add_57913_comb;
    p2_add_57914 <= p2_add_57914_comb;
    p2_add_57915 <= p2_add_57915_comb;
    p2_add_57916 <= p2_add_57916_comb;
    p2_add_57909 <= p2_add_57909_comb;
    p2_add_57910 <= p2_add_57910_comb;
    p2_add_57911 <= p2_add_57911_comb;
    p2_add_57912 <= p2_add_57912_comb;
    p2_add_57905 <= p2_add_57905_comb;
    p2_add_57906 <= p2_add_57906_comb;
    p2_add_57907 <= p2_add_57907_comb;
    p2_add_57908 <= p2_add_57908_comb;
    p2_add_57901 <= p2_add_57901_comb;
    p2_add_57902 <= p2_add_57902_comb;
    p2_add_57903 <= p2_add_57903_comb;
    p2_add_57904 <= p2_add_57904_comb;
    p2_add_57897 <= p2_add_57897_comb;
    p2_add_57898 <= p2_add_57898_comb;
    p2_add_57899 <= p2_add_57899_comb;
    p2_add_57900 <= p2_add_57900_comb;
    p2_add_57893 <= p2_add_57893_comb;
    p2_add_57894 <= p2_add_57894_comb;
    p2_add_57895 <= p2_add_57895_comb;
    p2_add_57896 <= p2_add_57896_comb;
    p2_add_57889 <= p2_add_57889_comb;
    p2_add_57890 <= p2_add_57890_comb;
    p2_add_57891 <= p2_add_57891_comb;
    p2_add_57892 <= p2_add_57892_comb;
    p2_add_57885 <= p2_add_57885_comb;
    p2_add_57886 <= p2_add_57886_comb;
    p2_add_57887 <= p2_add_57887_comb;
    p2_add_57888 <= p2_add_57888_comb;
    p2_add_57881 <= p2_add_57881_comb;
    p2_add_57882 <= p2_add_57882_comb;
    p2_add_57883 <= p2_add_57883_comb;
    p2_add_57884 <= p2_add_57884_comb;
    p2_add_57877 <= p2_add_57877_comb;
    p2_add_57878 <= p2_add_57878_comb;
    p2_add_57879 <= p2_add_57879_comb;
    p2_add_57880 <= p2_add_57880_comb;
    p2_add_57873 <= p2_add_57873_comb;
    p2_add_57874 <= p2_add_57874_comb;
    p2_add_57875 <= p2_add_57875_comb;
    p2_add_57876 <= p2_add_57876_comb;
    p2_add_57869 <= p2_add_57869_comb;
    p2_add_57870 <= p2_add_57870_comb;
    p2_add_57871 <= p2_add_57871_comb;
    p2_add_57872 <= p2_add_57872_comb;
    p2_add_57865 <= p2_add_57865_comb;
    p2_add_57866 <= p2_add_57866_comb;
    p2_add_57867 <= p2_add_57867_comb;
    p2_add_57868 <= p2_add_57868_comb;
    p2_add_57861 <= p2_add_57861_comb;
    p2_add_57862 <= p2_add_57862_comb;
    p2_add_57863 <= p2_add_57863_comb;
    p2_add_57864 <= p2_add_57864_comb;
    p2_add_57857 <= p2_add_57857_comb;
    p2_add_57858 <= p2_add_57858_comb;
    p2_add_57859 <= p2_add_57859_comb;
    p2_add_57860 <= p2_add_57860_comb;
    p2_add_57853 <= p2_add_57853_comb;
    p2_add_57854 <= p2_add_57854_comb;
    p2_add_57855 <= p2_add_57855_comb;
    p2_add_57856 <= p2_add_57856_comb;
    p2_add_57849 <= p2_add_57849_comb;
    p2_add_57850 <= p2_add_57850_comb;
    p2_add_57851 <= p2_add_57851_comb;
    p2_add_57852 <= p2_add_57852_comb;
  end

  // ===== Pipe stage 3:
  wire [31:0] p3_add_58621_comb;
  wire [31:0] p3_add_58622_comb;
  wire [31:0] p3_add_58623_comb;
  wire [31:0] p3_add_58624_comb;
  wire [31:0] p3_add_58625_comb;
  wire [31:0] p3_add_58626_comb;
  wire [31:0] p3_add_58627_comb;
  wire [31:0] p3_add_58628_comb;
  wire [31:0] p3_add_58629_comb;
  wire [31:0] p3_add_58630_comb;
  wire [31:0] p3_add_58631_comb;
  wire [31:0] p3_add_58632_comb;
  wire [31:0] p3_add_58633_comb;
  wire [31:0] p3_add_58634_comb;
  wire [31:0] p3_add_58635_comb;
  wire [31:0] p3_add_58636_comb;
  wire [31:0] p3_add_58637_comb;
  wire [31:0] p3_add_58638_comb;
  wire [31:0] p3_add_58639_comb;
  wire [31:0] p3_add_58640_comb;
  wire [31:0] p3_add_58641_comb;
  wire [31:0] p3_add_58642_comb;
  wire [31:0] p3_add_58643_comb;
  wire [31:0] p3_add_58644_comb;
  wire [31:0] p3_add_58645_comb;
  wire [31:0] p3_add_58646_comb;
  wire [31:0] p3_add_58647_comb;
  wire [31:0] p3_add_58648_comb;
  wire [31:0] p3_add_58649_comb;
  wire [31:0] p3_add_58650_comb;
  wire [31:0] p3_add_58651_comb;
  wire [31:0] p3_add_58652_comb;
  wire [31:0] p3_add_58653_comb;
  wire [31:0] p3_add_58654_comb;
  wire [31:0] p3_add_58655_comb;
  wire [31:0] p3_add_58656_comb;
  wire [31:0] p3_add_58657_comb;
  wire [31:0] p3_add_58658_comb;
  wire [31:0] p3_add_58659_comb;
  wire [31:0] p3_add_58660_comb;
  wire [31:0] p3_add_58661_comb;
  wire [31:0] p3_add_58662_comb;
  wire [31:0] p3_add_58663_comb;
  wire [31:0] p3_add_58664_comb;
  wire [31:0] p3_add_58665_comb;
  wire [31:0] p3_add_58666_comb;
  wire [31:0] p3_add_58667_comb;
  wire [31:0] p3_add_58668_comb;
  wire [31:0] p3_add_58669_comb;
  wire [31:0] p3_add_58670_comb;
  wire [31:0] p3_add_58671_comb;
  wire [31:0] p3_add_58672_comb;
  wire [31:0] p3_add_58673_comb;
  wire [31:0] p3_add_58674_comb;
  wire [31:0] p3_add_58675_comb;
  wire [31:0] p3_add_58676_comb;
  wire [31:0] p3_add_58677_comb;
  wire [31:0] p3_add_58678_comb;
  wire [31:0] p3_add_58679_comb;
  wire [31:0] p3_add_58680_comb;
  wire [31:0] p3_add_58681_comb;
  wire [31:0] p3_add_58682_comb;
  wire [31:0] p3_add_58683_comb;
  wire [31:0] p3_add_58684_comb;
  wire [31:0] p3_add_58685_comb;
  wire [31:0] p3_add_58686_comb;
  wire [31:0] p3_add_58687_comb;
  wire [31:0] p3_add_58688_comb;
  wire [31:0] p3_add_58689_comb;
  wire [31:0] p3_add_58690_comb;
  wire [31:0] p3_add_58691_comb;
  wire [31:0] p3_add_58692_comb;
  wire [31:0] p3_add_58693_comb;
  wire [31:0] p3_add_58694_comb;
  wire [31:0] p3_add_58695_comb;
  wire [31:0] p3_add_58696_comb;
  wire [31:0] p3_add_58697_comb;
  wire [31:0] p3_add_58698_comb;
  wire [31:0] p3_add_58699_comb;
  wire [31:0] p3_add_58700_comb;
  wire [31:0] p3_add_58701_comb;
  wire [31:0] p3_add_58702_comb;
  wire [31:0] p3_add_58703_comb;
  wire [31:0] p3_add_58704_comb;
  wire [31:0] p3_add_58705_comb;
  wire [31:0] p3_add_58706_comb;
  wire [31:0] p3_add_58707_comb;
  wire [31:0] p3_add_58708_comb;
  wire [31:0] p3_add_58709_comb;
  wire [31:0] p3_add_58710_comb;
  wire [31:0] p3_add_58711_comb;
  wire [31:0] p3_add_58712_comb;
  wire [31:0] p3_add_58713_comb;
  wire [31:0] p3_add_58714_comb;
  wire [31:0] p3_add_58715_comb;
  wire [31:0] p3_add_58716_comb;
  wire [31:0] p3_add_58717_comb;
  wire [31:0] p3_add_58718_comb;
  wire [31:0] p3_add_58719_comb;
  wire [31:0] p3_add_58720_comb;
  wire [31:0] p3_add_58721_comb;
  wire [31:0] p3_add_58722_comb;
  wire [31:0] p3_add_58723_comb;
  wire [31:0] p3_add_58724_comb;
  wire [31:0] p3_add_58725_comb;
  wire [31:0] p3_add_58726_comb;
  wire [31:0] p3_add_58727_comb;
  wire [31:0] p3_add_58728_comb;
  wire [31:0] p3_add_58729_comb;
  wire [31:0] p3_add_58730_comb;
  wire [31:0] p3_add_58731_comb;
  wire [31:0] p3_add_58732_comb;
  wire [31:0] p3_add_58733_comb;
  wire [31:0] p3_add_58734_comb;
  wire [31:0] p3_add_58735_comb;
  wire [31:0] p3_add_58736_comb;
  wire [31:0] p3_add_58737_comb;
  wire [31:0] p3_add_58738_comb;
  wire [31:0] p3_add_58739_comb;
  wire [31:0] p3_add_58740_comb;
  wire [31:0] p3_add_58741_comb;
  wire [31:0] p3_add_58742_comb;
  wire [31:0] p3_add_58743_comb;
  wire [31:0] p3_add_58744_comb;
  wire [31:0] p3_add_58745_comb;
  wire [31:0] p3_add_58746_comb;
  wire [31:0] p3_add_58747_comb;
  wire [31:0] p3_add_58748_comb;
  wire [31:0] p3_add_58749_comb;
  wire [31:0] p3_add_58750_comb;
  wire [31:0] p3_add_58751_comb;
  wire [31:0] p3_add_58752_comb;
  wire [31:0] p3_add_58753_comb;
  wire [31:0] p3_add_58754_comb;
  wire [31:0] p3_add_58755_comb;
  wire [31:0] p3_add_58756_comb;
  wire [31:0] p3_add_58757_comb;
  wire [31:0] p3_add_58758_comb;
  wire [31:0] p3_add_58759_comb;
  wire [31:0] p3_add_58760_comb;
  wire [31:0] p3_add_58761_comb;
  wire [31:0] p3_add_58762_comb;
  wire [31:0] p3_add_58763_comb;
  wire [31:0] p3_add_58764_comb;
  wire [31:0] p3_add_58765_comb;
  wire [31:0] p3_add_58766_comb;
  wire [31:0] p3_add_58767_comb;
  wire [31:0] p3_add_58768_comb;
  wire [31:0] p3_add_58769_comb;
  wire [31:0] p3_add_58770_comb;
  wire [31:0] p3_add_58771_comb;
  wire [31:0] p3_add_58772_comb;
  wire [31:0] p3_add_58773_comb;
  wire [31:0] p3_add_58774_comb;
  wire [31:0] p3_add_58775_comb;
  wire [31:0] p3_add_58776_comb;
  wire [31:0] p3_add_58777_comb;
  wire [31:0] p3_add_58778_comb;
  wire [31:0] p3_add_58779_comb;
  wire [31:0] p3_add_58780_comb;
  wire [31:0] p3_add_58781_comb;
  wire [31:0] p3_add_58782_comb;
  wire [31:0] p3_add_58783_comb;
  wire [31:0] p3_add_58784_comb;
  wire [31:0] p3_add_58785_comb;
  wire [31:0] p3_add_58786_comb;
  wire [31:0] p3_add_58787_comb;
  wire [31:0] p3_add_58788_comb;
  wire [31:0] p3_add_58789_comb;
  wire [31:0] p3_add_58790_comb;
  wire [31:0] p3_add_58791_comb;
  wire [31:0] p3_add_58792_comb;
  wire [31:0] p3_add_58793_comb;
  wire [31:0] p3_add_58794_comb;
  wire [31:0] p3_add_58795_comb;
  wire [31:0] p3_add_58796_comb;
  wire [31:0] p3_add_58797_comb;
  wire [31:0] p3_add_58798_comb;
  wire [31:0] p3_add_58799_comb;
  wire [31:0] p3_add_58800_comb;
  wire [31:0] p3_add_58801_comb;
  wire [31:0] p3_add_58802_comb;
  wire [31:0] p3_add_58803_comb;
  wire [31:0] p3_add_58804_comb;
  wire [31:0] p3_add_58805_comb;
  wire [31:0] p3_add_58806_comb;
  wire [31:0] p3_add_58807_comb;
  wire [31:0] p3_add_58808_comb;
  wire [31:0] p3_add_58809_comb;
  wire [31:0] p3_add_58810_comb;
  wire [31:0] p3_add_58811_comb;
  wire [31:0] p3_add_58812_comb;
  wire [31:0] p3_array_58813_comb[8];
  wire [31:0] p3_array_58814_comb[8];
  wire [31:0] p3_array_58815_comb[8];
  wire [31:0] p3_array_58816_comb[8];
  wire [31:0] p3_array_58817_comb[8];
  wire [31:0] p3_array_58818_comb[8];
  wire [31:0] p3_array_58819_comb[8];
  wire [31:0] p3_array_58820_comb[8];
  wire [31:0] p3_array_58821_comb[8][8];
  wire [6143:0] p3_tuple_58822_comb;
  assign p3_add_58621_comb = p2_add_57849 + p2_add_57850;
  assign p3_add_58622_comb = p2_add_57851 + p2_add_57852;
  assign p3_add_58623_comb = p2_add_57853 + p2_add_57854;
  assign p3_add_58624_comb = p2_add_57855 + p2_add_57856;
  assign p3_add_58625_comb = p2_add_57857 + p2_add_57858;
  assign p3_add_58626_comb = p2_add_57859 + p2_add_57860;
  assign p3_add_58627_comb = p2_add_57861 + p2_add_57862;
  assign p3_add_58628_comb = p2_add_57863 + p2_add_57864;
  assign p3_add_58629_comb = p2_add_57865 + p2_add_57866;
  assign p3_add_58630_comb = p2_add_57867 + p2_add_57868;
  assign p3_add_58631_comb = p2_add_57869 + p2_add_57870;
  assign p3_add_58632_comb = p2_add_57871 + p2_add_57872;
  assign p3_add_58633_comb = p2_add_57873 + p2_add_57874;
  assign p3_add_58634_comb = p2_add_57875 + p2_add_57876;
  assign p3_add_58635_comb = p2_add_57877 + p2_add_57878;
  assign p3_add_58636_comb = p2_add_57879 + p2_add_57880;
  assign p3_add_58637_comb = p2_add_57881 + p2_add_57882;
  assign p3_add_58638_comb = p2_add_57883 + p2_add_57884;
  assign p3_add_58639_comb = p2_add_57885 + p2_add_57886;
  assign p3_add_58640_comb = p2_add_57887 + p2_add_57888;
  assign p3_add_58641_comb = p2_add_57889 + p2_add_57890;
  assign p3_add_58642_comb = p2_add_57891 + p2_add_57892;
  assign p3_add_58643_comb = p2_add_57893 + p2_add_57894;
  assign p3_add_58644_comb = p2_add_57895 + p2_add_57896;
  assign p3_add_58645_comb = p2_add_57897 + p2_add_57898;
  assign p3_add_58646_comb = p2_add_57899 + p2_add_57900;
  assign p3_add_58647_comb = p2_add_57901 + p2_add_57902;
  assign p3_add_58648_comb = p2_add_57903 + p2_add_57904;
  assign p3_add_58649_comb = p2_add_57905 + p2_add_57906;
  assign p3_add_58650_comb = p2_add_57907 + p2_add_57908;
  assign p3_add_58651_comb = p2_add_57909 + p2_add_57910;
  assign p3_add_58652_comb = p2_add_57911 + p2_add_57912;
  assign p3_add_58653_comb = p2_add_57913 + p2_add_57914;
  assign p3_add_58654_comb = p2_add_57915 + p2_add_57916;
  assign p3_add_58655_comb = p2_add_57917 + p2_add_57918;
  assign p3_add_58656_comb = p2_add_57919 + p2_add_57920;
  assign p3_add_58657_comb = p2_add_57921 + p2_add_57922;
  assign p3_add_58658_comb = p2_add_57923 + p2_add_57924;
  assign p3_add_58659_comb = p2_add_57925 + p2_add_57926;
  assign p3_add_58660_comb = p2_add_57927 + p2_add_57928;
  assign p3_add_58661_comb = p2_add_57929 + p2_add_57930;
  assign p3_add_58662_comb = p2_add_57931 + p2_add_57932;
  assign p3_add_58663_comb = p2_add_57933 + p2_add_57934;
  assign p3_add_58664_comb = p2_add_57935 + p2_add_57936;
  assign p3_add_58665_comb = p2_add_57937 + p2_add_57938;
  assign p3_add_58666_comb = p2_add_57939 + p2_add_57940;
  assign p3_add_58667_comb = p2_add_57941 + p2_add_57942;
  assign p3_add_58668_comb = p2_add_57943 + p2_add_57944;
  assign p3_add_58669_comb = p2_add_57945 + p2_add_57946;
  assign p3_add_58670_comb = p2_add_57947 + p2_add_57948;
  assign p3_add_58671_comb = p2_add_57949 + p2_add_57950;
  assign p3_add_58672_comb = p2_add_57951 + p2_add_57952;
  assign p3_add_58673_comb = p2_add_57953 + p2_add_57954;
  assign p3_add_58674_comb = p2_add_57955 + p2_add_57956;
  assign p3_add_58675_comb = p2_add_57957 + p2_add_57958;
  assign p3_add_58676_comb = p2_add_57959 + p2_add_57960;
  assign p3_add_58677_comb = p2_add_57961 + p2_add_57962;
  assign p3_add_58678_comb = p2_add_57963 + p2_add_57964;
  assign p3_add_58679_comb = p2_add_57965 + p2_add_57966;
  assign p3_add_58680_comb = p2_add_57967 + p2_add_57968;
  assign p3_add_58681_comb = p2_add_57969 + p2_add_57970;
  assign p3_add_58682_comb = p2_add_57971 + p2_add_57972;
  assign p3_add_58683_comb = p2_add_57973 + p2_add_57974;
  assign p3_add_58684_comb = p2_add_57975 + p2_add_57976;
  assign p3_add_58685_comb = p2_add_57977 + p2_add_57978;
  assign p3_add_58686_comb = p2_add_57979 + p2_add_57980;
  assign p3_add_58687_comb = p2_add_57981 + p2_add_57982;
  assign p3_add_58688_comb = p2_add_57983 + p2_add_57984;
  assign p3_add_58689_comb = p2_add_57985 + p2_add_57986;
  assign p3_add_58690_comb = p2_add_57987 + p2_add_57988;
  assign p3_add_58691_comb = p2_add_57989 + p2_add_57990;
  assign p3_add_58692_comb = p2_add_57991 + p2_add_57992;
  assign p3_add_58693_comb = p2_add_57993 + p2_add_57994;
  assign p3_add_58694_comb = p2_add_57995 + p2_add_57996;
  assign p3_add_58695_comb = p2_add_57997 + p2_add_57998;
  assign p3_add_58696_comb = p2_add_57999 + p2_add_58000;
  assign p3_add_58697_comb = p2_add_58001 + p2_add_58002;
  assign p3_add_58698_comb = p2_add_58003 + p2_add_58004;
  assign p3_add_58699_comb = p2_add_58005 + p2_add_58006;
  assign p3_add_58700_comb = p2_add_58007 + p2_add_58008;
  assign p3_add_58701_comb = p2_add_58009 + p2_add_58010;
  assign p3_add_58702_comb = p2_add_58011 + p2_add_58012;
  assign p3_add_58703_comb = p2_add_58013 + p2_add_58014;
  assign p3_add_58704_comb = p2_add_58015 + p2_add_58016;
  assign p3_add_58705_comb = p2_add_58017 + p2_add_58018;
  assign p3_add_58706_comb = p2_add_58019 + p2_add_58020;
  assign p3_add_58707_comb = p2_add_58021 + p2_add_58022;
  assign p3_add_58708_comb = p2_add_58023 + p2_add_58024;
  assign p3_add_58709_comb = p2_add_58025 + p2_add_58026;
  assign p3_add_58710_comb = p2_add_58027 + p2_add_58028;
  assign p3_add_58711_comb = p2_add_58029 + p2_add_58030;
  assign p3_add_58712_comb = p2_add_58031 + p2_add_58032;
  assign p3_add_58713_comb = p2_add_58033 + p2_add_58034;
  assign p3_add_58714_comb = p2_add_58035 + p2_add_58036;
  assign p3_add_58715_comb = p2_add_58037 + p2_add_58038;
  assign p3_add_58716_comb = p2_add_58039 + p2_add_58040;
  assign p3_add_58717_comb = p2_add_58041 + p2_add_58042;
  assign p3_add_58718_comb = p2_add_58043 + p2_add_58044;
  assign p3_add_58719_comb = p2_add_58045 + p2_add_58046;
  assign p3_add_58720_comb = p2_add_58047 + p2_add_58048;
  assign p3_add_58721_comb = p2_add_58049 + p2_add_58050;
  assign p3_add_58722_comb = p2_add_58051 + p2_add_58052;
  assign p3_add_58723_comb = p2_add_58053 + p2_add_58054;
  assign p3_add_58724_comb = p2_add_58055 + p2_add_58056;
  assign p3_add_58725_comb = p2_add_58057 + p2_add_58058;
  assign p3_add_58726_comb = p2_add_58059 + p2_add_58060;
  assign p3_add_58727_comb = p2_add_58061 + p2_add_58062;
  assign p3_add_58728_comb = p2_add_58063 + p2_add_58064;
  assign p3_add_58729_comb = p2_add_58065 + p2_add_58066;
  assign p3_add_58730_comb = p2_add_58067 + p2_add_58068;
  assign p3_add_58731_comb = p2_add_58069 + p2_add_58070;
  assign p3_add_58732_comb = p2_add_58071 + p2_add_58072;
  assign p3_add_58733_comb = p2_add_58073 + p2_add_58074;
  assign p3_add_58734_comb = p2_add_58075 + p2_add_58076;
  assign p3_add_58735_comb = p2_add_58077 + p2_add_58078;
  assign p3_add_58736_comb = p2_add_58079 + p2_add_58080;
  assign p3_add_58737_comb = p2_add_58081 + p2_add_58082;
  assign p3_add_58738_comb = p2_add_58083 + p2_add_58084;
  assign p3_add_58739_comb = p2_add_58085 + p2_add_58086;
  assign p3_add_58740_comb = p2_add_58087 + p2_add_58088;
  assign p3_add_58741_comb = p2_add_58089 + p2_add_58090;
  assign p3_add_58742_comb = p2_add_58091 + p2_add_58092;
  assign p3_add_58743_comb = p2_add_58093 + p2_add_58094;
  assign p3_add_58744_comb = p2_add_58095 + p2_add_58096;
  assign p3_add_58745_comb = p2_add_58097 + p2_add_58098;
  assign p3_add_58746_comb = p2_add_58099 + p2_add_58100;
  assign p3_add_58747_comb = p2_add_58101 + p2_add_58102;
  assign p3_add_58748_comb = p2_add_58103 + p2_add_58104;
  assign p3_add_58749_comb = p3_add_58621_comb + p3_add_58622_comb;
  assign p3_add_58750_comb = p3_add_58623_comb + p3_add_58624_comb;
  assign p3_add_58751_comb = p3_add_58625_comb + p3_add_58626_comb;
  assign p3_add_58752_comb = p3_add_58627_comb + p3_add_58628_comb;
  assign p3_add_58753_comb = p3_add_58629_comb + p3_add_58630_comb;
  assign p3_add_58754_comb = p3_add_58631_comb + p3_add_58632_comb;
  assign p3_add_58755_comb = p3_add_58633_comb + p3_add_58634_comb;
  assign p3_add_58756_comb = p3_add_58635_comb + p3_add_58636_comb;
  assign p3_add_58757_comb = p3_add_58637_comb + p3_add_58638_comb;
  assign p3_add_58758_comb = p3_add_58639_comb + p3_add_58640_comb;
  assign p3_add_58759_comb = p3_add_58641_comb + p3_add_58642_comb;
  assign p3_add_58760_comb = p3_add_58643_comb + p3_add_58644_comb;
  assign p3_add_58761_comb = p3_add_58645_comb + p3_add_58646_comb;
  assign p3_add_58762_comb = p3_add_58647_comb + p3_add_58648_comb;
  assign p3_add_58763_comb = p3_add_58649_comb + p3_add_58650_comb;
  assign p3_add_58764_comb = p3_add_58651_comb + p3_add_58652_comb;
  assign p3_add_58765_comb = p3_add_58653_comb + p3_add_58654_comb;
  assign p3_add_58766_comb = p3_add_58655_comb + p3_add_58656_comb;
  assign p3_add_58767_comb = p3_add_58657_comb + p3_add_58658_comb;
  assign p3_add_58768_comb = p3_add_58659_comb + p3_add_58660_comb;
  assign p3_add_58769_comb = p3_add_58661_comb + p3_add_58662_comb;
  assign p3_add_58770_comb = p3_add_58663_comb + p3_add_58664_comb;
  assign p3_add_58771_comb = p3_add_58665_comb + p3_add_58666_comb;
  assign p3_add_58772_comb = p3_add_58667_comb + p3_add_58668_comb;
  assign p3_add_58773_comb = p3_add_58669_comb + p3_add_58670_comb;
  assign p3_add_58774_comb = p3_add_58671_comb + p3_add_58672_comb;
  assign p3_add_58775_comb = p3_add_58673_comb + p3_add_58674_comb;
  assign p3_add_58776_comb = p3_add_58675_comb + p3_add_58676_comb;
  assign p3_add_58777_comb = p3_add_58677_comb + p3_add_58678_comb;
  assign p3_add_58778_comb = p3_add_58679_comb + p3_add_58680_comb;
  assign p3_add_58779_comb = p3_add_58681_comb + p3_add_58682_comb;
  assign p3_add_58780_comb = p3_add_58683_comb + p3_add_58684_comb;
  assign p3_add_58781_comb = p3_add_58685_comb + p3_add_58686_comb;
  assign p3_add_58782_comb = p3_add_58687_comb + p3_add_58688_comb;
  assign p3_add_58783_comb = p3_add_58689_comb + p3_add_58690_comb;
  assign p3_add_58784_comb = p3_add_58691_comb + p3_add_58692_comb;
  assign p3_add_58785_comb = p3_add_58693_comb + p3_add_58694_comb;
  assign p3_add_58786_comb = p3_add_58695_comb + p3_add_58696_comb;
  assign p3_add_58787_comb = p3_add_58697_comb + p3_add_58698_comb;
  assign p3_add_58788_comb = p3_add_58699_comb + p3_add_58700_comb;
  assign p3_add_58789_comb = p3_add_58701_comb + p3_add_58702_comb;
  assign p3_add_58790_comb = p3_add_58703_comb + p3_add_58704_comb;
  assign p3_add_58791_comb = p3_add_58705_comb + p3_add_58706_comb;
  assign p3_add_58792_comb = p3_add_58707_comb + p3_add_58708_comb;
  assign p3_add_58793_comb = p3_add_58709_comb + p3_add_58710_comb;
  assign p3_add_58794_comb = p3_add_58711_comb + p3_add_58712_comb;
  assign p3_add_58795_comb = p3_add_58713_comb + p3_add_58714_comb;
  assign p3_add_58796_comb = p3_add_58715_comb + p3_add_58716_comb;
  assign p3_add_58797_comb = p3_add_58717_comb + p3_add_58718_comb;
  assign p3_add_58798_comb = p3_add_58719_comb + p3_add_58720_comb;
  assign p3_add_58799_comb = p3_add_58721_comb + p3_add_58722_comb;
  assign p3_add_58800_comb = p3_add_58723_comb + p3_add_58724_comb;
  assign p3_add_58801_comb = p3_add_58725_comb + p3_add_58726_comb;
  assign p3_add_58802_comb = p3_add_58727_comb + p3_add_58728_comb;
  assign p3_add_58803_comb = p3_add_58729_comb + p3_add_58730_comb;
  assign p3_add_58804_comb = p3_add_58731_comb + p3_add_58732_comb;
  assign p3_add_58805_comb = p3_add_58733_comb + p3_add_58734_comb;
  assign p3_add_58806_comb = p3_add_58735_comb + p3_add_58736_comb;
  assign p3_add_58807_comb = p3_add_58737_comb + p3_add_58738_comb;
  assign p3_add_58808_comb = p3_add_58739_comb + p3_add_58740_comb;
  assign p3_add_58809_comb = p3_add_58741_comb + p3_add_58742_comb;
  assign p3_add_58810_comb = p3_add_58743_comb + p3_add_58744_comb;
  assign p3_add_58811_comb = p3_add_58745_comb + p3_add_58746_comb;
  assign p3_add_58812_comb = p3_add_58747_comb + p3_add_58748_comb;
  assign p3_array_58813_comb[0] = p3_add_58749_comb;
  assign p3_array_58813_comb[1] = p3_add_58750_comb;
  assign p3_array_58813_comb[2] = p3_add_58751_comb;
  assign p3_array_58813_comb[3] = p3_add_58752_comb;
  assign p3_array_58813_comb[4] = p3_add_58753_comb;
  assign p3_array_58813_comb[5] = p3_add_58754_comb;
  assign p3_array_58813_comb[6] = p3_add_58755_comb;
  assign p3_array_58813_comb[7] = p3_add_58756_comb;
  assign p3_array_58814_comb[0] = p3_add_58757_comb;
  assign p3_array_58814_comb[1] = p3_add_58758_comb;
  assign p3_array_58814_comb[2] = p3_add_58759_comb;
  assign p3_array_58814_comb[3] = p3_add_58760_comb;
  assign p3_array_58814_comb[4] = p3_add_58761_comb;
  assign p3_array_58814_comb[5] = p3_add_58762_comb;
  assign p3_array_58814_comb[6] = p3_add_58763_comb;
  assign p3_array_58814_comb[7] = p3_add_58764_comb;
  assign p3_array_58815_comb[0] = p3_add_58765_comb;
  assign p3_array_58815_comb[1] = p3_add_58766_comb;
  assign p3_array_58815_comb[2] = p3_add_58767_comb;
  assign p3_array_58815_comb[3] = p3_add_58768_comb;
  assign p3_array_58815_comb[4] = p3_add_58769_comb;
  assign p3_array_58815_comb[5] = p3_add_58770_comb;
  assign p3_array_58815_comb[6] = p3_add_58771_comb;
  assign p3_array_58815_comb[7] = p3_add_58772_comb;
  assign p3_array_58816_comb[0] = p3_add_58773_comb;
  assign p3_array_58816_comb[1] = p3_add_58774_comb;
  assign p3_array_58816_comb[2] = p3_add_58775_comb;
  assign p3_array_58816_comb[3] = p3_add_58776_comb;
  assign p3_array_58816_comb[4] = p3_add_58777_comb;
  assign p3_array_58816_comb[5] = p3_add_58778_comb;
  assign p3_array_58816_comb[6] = p3_add_58779_comb;
  assign p3_array_58816_comb[7] = p3_add_58780_comb;
  assign p3_array_58817_comb[0] = p3_add_58781_comb;
  assign p3_array_58817_comb[1] = p3_add_58782_comb;
  assign p3_array_58817_comb[2] = p3_add_58783_comb;
  assign p3_array_58817_comb[3] = p3_add_58784_comb;
  assign p3_array_58817_comb[4] = p3_add_58785_comb;
  assign p3_array_58817_comb[5] = p3_add_58786_comb;
  assign p3_array_58817_comb[6] = p3_add_58787_comb;
  assign p3_array_58817_comb[7] = p3_add_58788_comb;
  assign p3_array_58818_comb[0] = p3_add_58789_comb;
  assign p3_array_58818_comb[1] = p3_add_58790_comb;
  assign p3_array_58818_comb[2] = p3_add_58791_comb;
  assign p3_array_58818_comb[3] = p3_add_58792_comb;
  assign p3_array_58818_comb[4] = p3_add_58793_comb;
  assign p3_array_58818_comb[5] = p3_add_58794_comb;
  assign p3_array_58818_comb[6] = p3_add_58795_comb;
  assign p3_array_58818_comb[7] = p3_add_58796_comb;
  assign p3_array_58819_comb[0] = p3_add_58797_comb;
  assign p3_array_58819_comb[1] = p3_add_58798_comb;
  assign p3_array_58819_comb[2] = p3_add_58799_comb;
  assign p3_array_58819_comb[3] = p3_add_58800_comb;
  assign p3_array_58819_comb[4] = p3_add_58801_comb;
  assign p3_array_58819_comb[5] = p3_add_58802_comb;
  assign p3_array_58819_comb[6] = p3_add_58803_comb;
  assign p3_array_58819_comb[7] = p3_add_58804_comb;
  assign p3_array_58820_comb[0] = p3_add_58805_comb;
  assign p3_array_58820_comb[1] = p3_add_58806_comb;
  assign p3_array_58820_comb[2] = p3_add_58807_comb;
  assign p3_array_58820_comb[3] = p3_add_58808_comb;
  assign p3_array_58820_comb[4] = p3_add_58809_comb;
  assign p3_array_58820_comb[5] = p3_add_58810_comb;
  assign p3_array_58820_comb[6] = p3_add_58811_comb;
  assign p3_array_58820_comb[7] = p3_add_58812_comb;
  assign p3_array_58821_comb[0] = p3_array_58813_comb;
  assign p3_array_58821_comb[1] = p3_array_58814_comb;
  assign p3_array_58821_comb[2] = p3_array_58815_comb;
  assign p3_array_58821_comb[3] = p3_array_58816_comb;
  assign p3_array_58821_comb[4] = p3_array_58817_comb;
  assign p3_array_58821_comb[5] = p3_array_58818_comb;
  assign p3_array_58821_comb[6] = p3_array_58819_comb;
  assign p3_array_58821_comb[7] = p3_array_58820_comb;
  assign p3_tuple_58822_comb = {{{p2_a[7][7], p2_a[7][6], p2_a[7][5], p2_a[7][4], p2_a[7][3], p2_a[7][2], p2_a[7][1], p2_a[7][0]}, {p2_a[6][7], p2_a[6][6], p2_a[6][5], p2_a[6][4], p2_a[6][3], p2_a[6][2], p2_a[6][1], p2_a[6][0]}, {p2_a[5][7], p2_a[5][6], p2_a[5][5], p2_a[5][4], p2_a[5][3], p2_a[5][2], p2_a[5][1], p2_a[5][0]}, {p2_a[4][7], p2_a[4][6], p2_a[4][5], p2_a[4][4], p2_a[4][3], p2_a[4][2], p2_a[4][1], p2_a[4][0]}, {p2_a[3][7], p2_a[3][6], p2_a[3][5], p2_a[3][4], p2_a[3][3], p2_a[3][2], p2_a[3][1], p2_a[3][0]}, {p2_a[2][7], p2_a[2][6], p2_a[2][5], p2_a[2][4], p2_a[2][3], p2_a[2][2], p2_a[2][1], p2_a[2][0]}, {p2_a[1][7], p2_a[1][6], p2_a[1][5], p2_a[1][4], p2_a[1][3], p2_a[1][2], p2_a[1][1], p2_a[1][0]}, {p2_a[0][7], p2_a[0][6], p2_a[0][5], p2_a[0][4], p2_a[0][3], p2_a[0][2], p2_a[0][1], p2_a[0][0]}}, {{p2_b[7][7], p2_b[7][6], p2_b[7][5], p2_b[7][4], p2_b[7][3], p2_b[7][2], p2_b[7][1], p2_b[7][0]}, {p2_b[6][7], p2_b[6][6], p2_b[6][5], p2_b[6][4], p2_b[6][3], p2_b[6][2], p2_b[6][1], p2_b[6][0]}, {p2_b[5][7], p2_b[5][6], p2_b[5][5], p2_b[5][4], p2_b[5][3], p2_b[5][2], p2_b[5][1], p2_b[5][0]}, {p2_b[4][7], p2_b[4][6], p2_b[4][5], p2_b[4][4], p2_b[4][3], p2_b[4][2], p2_b[4][1], p2_b[4][0]}, {p2_b[3][7], p2_b[3][6], p2_b[3][5], p2_b[3][4], p2_b[3][3], p2_b[3][2], p2_b[3][1], p2_b[3][0]}, {p2_b[2][7], p2_b[2][6], p2_b[2][5], p2_b[2][4], p2_b[2][3], p2_b[2][2], p2_b[2][1], p2_b[2][0]}, {p2_b[1][7], p2_b[1][6], p2_b[1][5], p2_b[1][4], p2_b[1][3], p2_b[1][2], p2_b[1][1], p2_b[1][0]}, {p2_b[0][7], p2_b[0][6], p2_b[0][5], p2_b[0][4], p2_b[0][3], p2_b[0][2], p2_b[0][1], p2_b[0][0]}}, {{p3_array_58821_comb[7][7], p3_array_58821_comb[7][6], p3_array_58821_comb[7][5], p3_array_58821_comb[7][4], p3_array_58821_comb[7][3], p3_array_58821_comb[7][2], p3_array_58821_comb[7][1], p3_array_58821_comb[7][0]}, {p3_array_58821_comb[6][7], p3_array_58821_comb[6][6], p3_array_58821_comb[6][5], p3_array_58821_comb[6][4], p3_array_58821_comb[6][3], p3_array_58821_comb[6][2], p3_array_58821_comb[6][1], p3_array_58821_comb[6][0]}, {p3_array_58821_comb[5][7], p3_array_58821_comb[5][6], p3_array_58821_comb[5][5], p3_array_58821_comb[5][4], p3_array_58821_comb[5][3], p3_array_58821_comb[5][2], p3_array_58821_comb[5][1], p3_array_58821_comb[5][0]}, {p3_array_58821_comb[4][7], p3_array_58821_comb[4][6], p3_array_58821_comb[4][5], p3_array_58821_comb[4][4], p3_array_58821_comb[4][3], p3_array_58821_comb[4][2], p3_array_58821_comb[4][1], p3_array_58821_comb[4][0]}, {p3_array_58821_comb[3][7], p3_array_58821_comb[3][6], p3_array_58821_comb[3][5], p3_array_58821_comb[3][4], p3_array_58821_comb[3][3], p3_array_58821_comb[3][2], p3_array_58821_comb[3][1], p3_array_58821_comb[3][0]}, {p3_array_58821_comb[2][7], p3_array_58821_comb[2][6], p3_array_58821_comb[2][5], p3_array_58821_comb[2][4], p3_array_58821_comb[2][3], p3_array_58821_comb[2][2], p3_array_58821_comb[2][1], p3_array_58821_comb[2][0]}, {p3_array_58821_comb[1][7], p3_array_58821_comb[1][6], p3_array_58821_comb[1][5], p3_array_58821_comb[1][4], p3_array_58821_comb[1][3], p3_array_58821_comb[1][2], p3_array_58821_comb[1][1], p3_array_58821_comb[1][0]}, {p3_array_58821_comb[0][7], p3_array_58821_comb[0][6], p3_array_58821_comb[0][5], p3_array_58821_comb[0][4], p3_array_58821_comb[0][3], p3_array_58821_comb[0][2], p3_array_58821_comb[0][1], p3_array_58821_comb[0][0]}}};

  // Registers for pipe stage 3:
  reg [6143:0] p3_tuple_58822;
  always_ff @ (posedge clk) begin
    p3_tuple_58822 <= p3_tuple_58822_comb;
  end
  assign out = p3_tuple_58822;
endmodule
