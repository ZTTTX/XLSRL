module xls_test(
  input wire clk,
  input wire [511:0] message,
  output wire [255:0] out
);
  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [511:0] p0_message;
  always_ff @ (posedge clk) begin
    p0_message <= message;
  end

  // ===== Pipe stage 1:
  wire [28:0] p1_add_62950_comb;
  wire [30:0] p1_add_62954_comb;
  wire [29:0] p1_add_62957_comb;
  assign p1_add_62950_comb = p0_message[511:483] + 29'h1e6e_fdad;
  assign p1_add_62954_comb = {p1_add_62950_comb, p0_message[482:481]} + 31'h52a7_fa9d;
  assign p1_add_62957_comb = p0_message[479:450] + 30'h242e_c78f;

  // Registers for pipe stage 1:
  reg [511:0] p1_message;
  reg [28:0] p1_add_62950;
  reg [30:0] p1_add_62954;
  reg [29:0] p1_add_62957;
  always_ff @ (posedge clk) begin
    p1_message <= p0_message;
    p1_add_62950 <= p1_add_62950_comb;
    p1_add_62954 <= p1_add_62954_comb;
    p1_add_62957 <= p1_add_62957_comb;
  end

  // ===== Pipe stage 2:
  wire p2_bit_slice_62966_comb;
  wire [31:0] p2_concat_62967_comb;
  wire [31:0] p2_add_62994_comb;
  wire [31:0] p2_add_62996_comb;
  wire [30:0] p2_add_62999_comb;
  assign p2_bit_slice_62966_comb = p1_message[480];
  assign p2_concat_62967_comb = {p1_add_62954, p2_bit_slice_62966_comb};
  assign p2_add_62994_comb = (p2_concat_62967_comb & 32'h510e_527f ^ ~(p2_concat_62967_comb | 32'h64fa_9773)) + {p1_add_62957, p1_message[449:448]};
  assign p2_add_62996_comb = p2_add_62994_comb + {{p1_add_62954[4:0], p2_bit_slice_62966_comb} ^ p1_add_62954[9:4] ^ p1_add_62954[23:18], p1_add_62954[30:26] ^ {p1_add_62954[3:0], p2_bit_slice_62966_comb} ^ p1_add_62954[17:13], p1_add_62954[25:12] ^ p1_add_62954[30:17] ^ {p1_add_62954[12:0], p2_bit_slice_62966_comb}, p1_add_62954[11:5] ^ p1_add_62954[16:10] ^ p1_add_62954[30:24]};
  assign p2_add_62999_comb = p2_add_62996_comb[31:1] + 31'h1e37_79b9;

  // Registers for pipe stage 2:
  reg [511:0] p2_message;
  reg p2_bit_slice_62966;
  reg [31:0] p2_concat_62967;
  reg [31:0] p2_add_62996;
  reg [28:0] p2_add_62950;
  reg [30:0] p2_add_62954;
  reg [30:0] p2_add_62999;
  always_ff @ (posedge clk) begin
    p2_message <= p1_message;
    p2_bit_slice_62966 <= p2_bit_slice_62966_comb;
    p2_concat_62967 <= p2_concat_62967_comb;
    p2_add_62996 <= p2_add_62996_comb;
    p2_add_62950 <= p1_add_62950;
    p2_add_62954 <= p1_add_62954;
    p2_add_62999 <= p2_add_62999_comb;
  end

  // ===== Pipe stage 3:
  wire [31:0] p3_concat_63020_comb;
  wire [31:0] p3_bit_slice_63040_comb;
  wire [31:0] p3_add_63062_comb;
  wire [31:0] p3_add_63044_comb;
  wire [31:0] p3_add_63045_comb;
  wire [31:0] p3_and_63065_comb;
  wire [31:0] p3_add_63046_comb;
  wire [31:0] p3_add_63050_comb;
  wire [31:0] p3_add_63085_comb;
  wire [31:0] p3_nor_63054_comb;
  wire [31:0] p3_concat_63058_comb;
  wire [31:0] p3_add_63087_comb;
  wire [29:0] p3_add_63055_comb;
  assign p3_concat_63020_comb = {p2_add_62999, p2_add_62996[0]};
  assign p3_bit_slice_63040_comb = p2_message[447:416];
  assign p3_add_63062_comb = {p2_add_62950, p2_message[482:480]} + 32'h0890_9ae5;
  assign p3_add_63044_comb = p3_bit_slice_63040_comb + ({p2_add_62999 & p2_add_62954, p2_add_62996[0] & p2_bit_slice_62966} ^ ~(p3_concat_63020_comb | 32'haef1_ad80));
  assign p3_add_63045_comb = {{p2_add_62999[4:0], p2_add_62996[0]} ^ p2_add_62999[9:4] ^ p2_add_62999[23:18], p2_add_62999[30:26] ^ {p2_add_62999[3:0], p2_add_62996[0]} ^ p2_add_62999[17:13], p2_add_62999[25:12] ^ p2_add_62999[30:17] ^ {p2_add_62999[12:0], p2_add_62996[0]}, p2_add_62999[11:5] ^ p2_add_62999[16:10] ^ p2_add_62999[30:24]} + 32'h50c6_645b;
  assign p3_and_63065_comb = p3_add_63062_comb & 32'h6a09_e667;
  assign p3_add_63046_comb = p3_add_63044_comb + p3_add_63045_comb;
  assign p3_add_63050_comb = p3_add_63046_comb + 32'hbb67_ae85;
  assign p3_add_63085_comb = (p3_and_63065_comb ^ p3_add_63062_comb & 32'hbb67_ae85 ^ 32'h2a01_a605) + p2_add_62996;
  assign p3_nor_63054_comb = ~(p3_add_63050_comb | {~p2_add_62954, ~p2_bit_slice_62966});
  assign p3_concat_63058_comb = {~p2_add_62999, ~p2_add_62996[0]};
  assign p3_add_63087_comb = p3_add_63085_comb + {p3_add_63062_comb[1:0] ^ p3_add_63062_comb[12:11] ^ p3_add_63062_comb[21:20], p3_add_63062_comb[31:21] ^ p3_add_63062_comb[10:0] ^ p3_add_63062_comb[19:9], p3_add_63062_comb[20:12] ^ p3_add_63062_comb[31:23] ^ p3_add_63062_comb[8:0], p3_add_63062_comb[11:2] ^ p3_add_63062_comb[22:13] ^ p3_add_63062_comb[31:22]};
  assign p3_add_63055_comb = p2_message[415:386] + 30'h0eb1_0b89;

  // Registers for pipe stage 3:
  reg [511:0] p3_message;
  reg [31:0] p3_concat_62967;
  reg [31:0] p3_concat_63020;
  reg [31:0] p3_bit_slice_63040;
  reg [31:0] p3_add_63046;
  reg [31:0] p3_nor_63054;
  reg [31:0] p3_concat_63058;
  reg [31:0] p3_and_63065;
  reg [31:0] p3_add_63087;
  reg [31:0] p3_add_63050;
  reg [29:0] p3_add_63055;
  reg [31:0] p3_add_63062;
  always_ff @ (posedge clk) begin
    p3_message <= p2_message;
    p3_concat_62967 <= p2_concat_62967;
    p3_concat_63020 <= p3_concat_63020_comb;
    p3_bit_slice_63040 <= p3_bit_slice_63040_comb;
    p3_add_63046 <= p3_add_63046_comb;
    p3_nor_63054 <= p3_nor_63054_comb;
    p3_concat_63058 <= p3_concat_63058_comb;
    p3_and_63065 <= p3_and_63065_comb;
    p3_add_63087 <= p3_add_63087_comb;
    p3_add_63050 <= p3_add_63050_comb;
    p3_add_63055 <= p3_add_63055_comb;
    p3_add_63062 <= p3_add_63062_comb;
  end

  // ===== Pipe stage 4:
  wire [31:0] p4_add_63132_comb;
  wire [31:0] p4_and_63143_comb;
  wire [31:0] p4_add_63134_comb;
  wire [31:0] p4_bit_slice_63138_comb;
  wire [31:0] p4_add_63136_comb;
  wire [31:0] p4_add_63140_comb;
  wire [31:0] p4_add_63162_comb;
  wire [31:0] p4_nor_63137_comb;
  wire [31:0] p4_add_63141_comb;
  wire [31:0] p4_add_63164_comb;
  assign p4_add_63132_comb = (p3_add_63050 & p3_concat_63020 ^ p3_nor_63054) + {p3_add_63055, p3_message[385:384]};
  assign p4_and_63143_comb = p3_add_63087 & p3_add_63062;
  assign p4_add_63134_comb = p4_add_63132_comb + {p3_add_63050[5:0] ^ p3_add_63050[10:5] ^ p3_add_63050[24:19], p3_add_63050[31:27] ^ p3_add_63050[4:0] ^ p3_add_63050[18:14], p3_add_63050[26:13] ^ p3_add_63050[31:18] ^ p3_add_63050[13:0], p3_add_63050[12:6] ^ p3_add_63050[17:11] ^ p3_add_63050[31:25]};
  assign p4_bit_slice_63138_comb = p3_message[383:352];
  assign p4_add_63136_comb = p4_add_63134_comb + 32'h6a09_e667;
  assign p4_add_63140_comb = p4_bit_slice_63138_comb + 32'h3956_c25b;
  assign p4_add_63162_comb = (p4_and_63143_comb ^ p3_add_63087 & 32'h6a09_e667 ^ p3_and_63065) + p3_add_63046;
  assign p4_nor_63137_comb = ~(p4_add_63136_comb | p3_concat_63058);
  assign p4_add_63141_comb = p3_concat_62967 + p4_add_63140_comb;
  assign p4_add_63164_comb = p4_add_63162_comb + {p3_add_63087[1:0] ^ p3_add_63087[12:11] ^ p3_add_63087[21:20], p3_add_63087[31:21] ^ p3_add_63087[10:0] ^ p3_add_63087[19:9], p3_add_63087[20:12] ^ p3_add_63087[31:23] ^ p3_add_63087[8:0], p3_add_63087[11:2] ^ p3_add_63087[22:13] ^ p3_add_63087[31:22]};

  // Registers for pipe stage 4:
  reg [511:0] p4_message;
  reg [31:0] p4_concat_63020;
  reg [31:0] p4_bit_slice_63040;
  reg [31:0] p4_add_63134;
  reg [31:0] p4_nor_63137;
  reg [31:0] p4_bit_slice_63138;
  reg [31:0] p4_add_63141;
  reg [31:0] p4_add_63087;
  reg [31:0] p4_and_63143;
  reg [31:0] p4_add_63164;
  reg [31:0] p4_add_63050;
  reg [31:0] p4_add_63136;
  reg [31:0] p4_add_63062;
  always_ff @ (posedge clk) begin
    p4_message <= p3_message;
    p4_concat_63020 <= p3_concat_63020;
    p4_bit_slice_63040 <= p3_bit_slice_63040;
    p4_add_63134 <= p4_add_63134_comb;
    p4_nor_63137 <= p4_nor_63137_comb;
    p4_bit_slice_63138 <= p4_bit_slice_63138_comb;
    p4_add_63141 <= p4_add_63141_comb;
    p4_add_63087 <= p3_add_63087;
    p4_and_63143 <= p4_and_63143_comb;
    p4_add_63164 <= p4_add_63164_comb;
    p4_add_63050 <= p3_add_63050;
    p4_add_63136 <= p4_add_63136_comb;
    p4_add_63062 <= p3_add_63062;
  end

  // ===== Pipe stage 5:
  wire [31:0] p5_and_63217_comb;
  wire [31:0] p5_add_63210_comb;
  wire [31:0] p5_bit_slice_63213_comb;
  wire [31:0] p5_add_63211_comb;
  wire [31:0] p5_add_63215_comb;
  wire [31:0] p5_add_63236_comb;
  wire [31:0] p5_add_63212_comb;
  wire [31:0] p5_add_63216_comb;
  wire [31:0] p5_add_63238_comb;
  assign p5_and_63217_comb = p4_add_63164 & p4_add_63087;
  assign p5_add_63210_comb = {p4_add_63136[5:0] ^ p4_add_63136[10:5] ^ p4_add_63136[24:19], p4_add_63136[31:27] ^ p4_add_63136[4:0] ^ p4_add_63136[18:14], p4_add_63136[26:13] ^ p4_add_63136[31:18] ^ p4_add_63136[13:0], p4_add_63136[12:6] ^ p4_add_63136[17:11] ^ p4_add_63136[31:25]} + (p4_add_63136 & p4_add_63050 ^ p4_nor_63137);
  assign p5_bit_slice_63213_comb = p4_message[351:320];
  assign p5_add_63211_comb = p5_add_63210_comb + p4_add_63141;
  assign p5_add_63215_comb = p5_bit_slice_63213_comb + 32'h59f1_11f1;
  assign p5_add_63236_comb = (p5_and_63217_comb ^ p4_add_63164 & p4_add_63062 ^ p4_and_63143) + p4_add_63134;
  assign p5_add_63212_comb = p5_add_63211_comb + p4_add_63062;
  assign p5_add_63216_comb = p4_concat_63020 + p5_add_63215_comb;
  assign p5_add_63238_comb = p5_add_63236_comb + {p4_add_63164[1:0] ^ p4_add_63164[12:11] ^ p4_add_63164[21:20], p4_add_63164[31:21] ^ p4_add_63164[10:0] ^ p4_add_63164[19:9], p4_add_63164[20:12] ^ p4_add_63164[31:23] ^ p4_add_63164[8:0], p4_add_63164[11:2] ^ p4_add_63164[22:13] ^ p4_add_63164[31:22]};

  // Registers for pipe stage 5:
  reg [511:0] p5_message;
  reg [31:0] p5_bit_slice_63040;
  reg [31:0] p5_bit_slice_63138;
  reg [31:0] p5_add_63211;
  reg [31:0] p5_add_63212;
  reg [31:0] p5_bit_slice_63213;
  reg [31:0] p5_add_63216;
  reg [31:0] p5_add_63087;
  reg [31:0] p5_add_63164;
  reg [31:0] p5_and_63217;
  reg [31:0] p5_add_63238;
  reg [31:0] p5_add_63050;
  reg [31:0] p5_add_63136;
  always_ff @ (posedge clk) begin
    p5_message <= p4_message;
    p5_bit_slice_63040 <= p4_bit_slice_63040;
    p5_bit_slice_63138 <= p4_bit_slice_63138;
    p5_add_63211 <= p5_add_63211_comb;
    p5_add_63212 <= p5_add_63212_comb;
    p5_bit_slice_63213 <= p5_bit_slice_63213_comb;
    p5_add_63216 <= p5_add_63216_comb;
    p5_add_63087 <= p4_add_63087;
    p5_add_63164 <= p4_add_63164;
    p5_and_63217 <= p5_and_63217_comb;
    p5_add_63238 <= p5_add_63238_comb;
    p5_add_63050 <= p4_add_63050;
    p5_add_63136 <= p4_add_63136;
  end

  // ===== Pipe stage 6:
  wire [31:0] p6_and_63295_comb;
  wire [31:0] p6_add_63286_comb;
  wire [29:0] p6_add_63291_comb;
  wire [31:0] p6_add_63287_comb;
  wire [31:0] p6_add_63314_comb;
  wire [31:0] p6_add_63288_comb;
  wire [31:0] p6_add_63294_comb;
  wire [31:0] p6_add_63316_comb;
  assign p6_and_63295_comb = p5_add_63238 & p5_add_63164;
  assign p6_add_63286_comb = {p5_add_63212[5:0] ^ p5_add_63212[10:5] ^ p5_add_63212[24:19], p5_add_63212[31:27] ^ p5_add_63212[4:0] ^ p5_add_63212[18:14], p5_add_63212[26:13] ^ p5_add_63212[31:18] ^ p5_add_63212[13:0], p5_add_63212[12:6] ^ p5_add_63212[17:11] ^ p5_add_63212[31:25]} + (p5_add_63212 & p5_add_63136 ^ ~(p5_add_63212 | ~p5_add_63050));
  assign p6_add_63291_comb = p5_message[319:290] + 30'h248f_e0a9;
  assign p6_add_63287_comb = p6_add_63286_comb + p5_add_63216;
  assign p6_add_63314_comb = (p6_and_63295_comb ^ p5_add_63238 & p5_add_63087 ^ p5_and_63217) + p5_add_63211;
  assign p6_add_63288_comb = p6_add_63287_comb + p5_add_63087;
  assign p6_add_63294_comb = {p6_add_63291_comb, p5_message[289:288]} + p5_add_63050;
  assign p6_add_63316_comb = p6_add_63314_comb + {p5_add_63238[1:0] ^ p5_add_63238[12:11] ^ p5_add_63238[21:20], p5_add_63238[31:21] ^ p5_add_63238[10:0] ^ p5_add_63238[19:9], p5_add_63238[20:12] ^ p5_add_63238[31:23] ^ p5_add_63238[8:0], p5_add_63238[11:2] ^ p5_add_63238[22:13] ^ p5_add_63238[31:22]};

  // Registers for pipe stage 6:
  reg [511:0] p6_message;
  reg [31:0] p6_bit_slice_63040;
  reg [31:0] p6_bit_slice_63138;
  reg [31:0] p6_add_63212;
  reg [31:0] p6_bit_slice_63213;
  reg [31:0] p6_add_63287;
  reg [31:0] p6_add_63288;
  reg [31:0] p6_add_63294;
  reg [31:0] p6_add_63164;
  reg [31:0] p6_add_63238;
  reg [31:0] p6_and_63295;
  reg [31:0] p6_add_63316;
  reg [31:0] p6_add_63136;
  always_ff @ (posedge clk) begin
    p6_message <= p5_message;
    p6_bit_slice_63040 <= p5_bit_slice_63040;
    p6_bit_slice_63138 <= p5_bit_slice_63138;
    p6_add_63212 <= p5_add_63212;
    p6_bit_slice_63213 <= p5_bit_slice_63213;
    p6_add_63287 <= p6_add_63287_comb;
    p6_add_63288 <= p6_add_63288_comb;
    p6_add_63294 <= p6_add_63294_comb;
    p6_add_63164 <= p5_add_63164;
    p6_add_63238 <= p5_add_63238;
    p6_and_63295 <= p6_and_63295_comb;
    p6_add_63316 <= p6_add_63316_comb;
    p6_add_63136 <= p5_add_63136;
  end

  // ===== Pipe stage 7:
  wire [31:0] p7_and_63371_comb;
  wire [31:0] p7_add_63364_comb;
  wire [31:0] p7_bit_slice_63367_comb;
  wire [31:0] p7_add_63365_comb;
  wire [31:0] p7_add_63369_comb;
  wire [31:0] p7_add_63390_comb;
  wire [31:0] p7_add_63366_comb;
  wire [31:0] p7_add_63370_comb;
  wire [31:0] p7_add_63392_comb;
  assign p7_and_63371_comb = p6_add_63316 & p6_add_63238;
  assign p7_add_63364_comb = (p6_add_63288 & p6_add_63212 ^ ~(p6_add_63288 | ~p6_add_63136)) + {p6_add_63288[5:0] ^ p6_add_63288[10:5] ^ p6_add_63288[24:19], p6_add_63288[31:27] ^ p6_add_63288[4:0] ^ p6_add_63288[18:14], p6_add_63288[26:13] ^ p6_add_63288[31:18] ^ p6_add_63288[13:0], p6_add_63288[12:6] ^ p6_add_63288[17:11] ^ p6_add_63288[31:25]};
  assign p7_bit_slice_63367_comb = p6_message[287:256];
  assign p7_add_63365_comb = p7_add_63364_comb + p6_add_63294;
  assign p7_add_63369_comb = p7_bit_slice_63367_comb + 32'hab1c_5ed5;
  assign p7_add_63390_comb = (p7_and_63371_comb ^ p6_add_63316 & p6_add_63164 ^ p6_and_63295) + p6_add_63287;
  assign p7_add_63366_comb = p7_add_63365_comb + p6_add_63164;
  assign p7_add_63370_comb = p6_add_63136 + p7_add_63369_comb;
  assign p7_add_63392_comb = p7_add_63390_comb + {p6_add_63316[1:0] ^ p6_add_63316[12:11] ^ p6_add_63316[21:20], p6_add_63316[31:21] ^ p6_add_63316[10:0] ^ p6_add_63316[19:9], p6_add_63316[20:12] ^ p6_add_63316[31:23] ^ p6_add_63316[8:0], p6_add_63316[11:2] ^ p6_add_63316[22:13] ^ p6_add_63316[31:22]};

  // Registers for pipe stage 7:
  reg [511:0] p7_message;
  reg [31:0] p7_bit_slice_63040;
  reg [31:0] p7_bit_slice_63138;
  reg [31:0] p7_add_63212;
  reg [31:0] p7_bit_slice_63213;
  reg [31:0] p7_add_63288;
  reg [31:0] p7_add_63365;
  reg [31:0] p7_add_63366;
  reg [31:0] p7_bit_slice_63367;
  reg [31:0] p7_add_63370;
  reg [31:0] p7_add_63238;
  reg [31:0] p7_add_63316;
  reg [31:0] p7_and_63371;
  reg [31:0] p7_add_63392;
  always_ff @ (posedge clk) begin
    p7_message <= p6_message;
    p7_bit_slice_63040 <= p6_bit_slice_63040;
    p7_bit_slice_63138 <= p6_bit_slice_63138;
    p7_add_63212 <= p6_add_63212;
    p7_bit_slice_63213 <= p6_bit_slice_63213;
    p7_add_63288 <= p6_add_63288;
    p7_add_63365 <= p7_add_63365_comb;
    p7_add_63366 <= p7_add_63366_comb;
    p7_bit_slice_63367 <= p7_bit_slice_63367_comb;
    p7_add_63370 <= p7_add_63370_comb;
    p7_add_63238 <= p6_add_63238;
    p7_add_63316 <= p6_add_63316;
    p7_and_63371 <= p7_and_63371_comb;
    p7_add_63392 <= p7_add_63392_comb;
  end

  // ===== Pipe stage 8:
  wire [31:0] p8_and_63451_comb;
  wire [31:0] p8_add_63442_comb;
  wire [28:0] p8_add_63447_comb;
  wire [31:0] p8_add_63443_comb;
  wire [31:0] p8_add_63470_comb;
  wire [31:0] p8_add_63444_comb;
  wire [31:0] p8_add_63450_comb;
  wire [31:0] p8_add_63472_comb;
  assign p8_and_63451_comb = p7_add_63392 & p7_add_63316;
  assign p8_add_63442_comb = {p7_add_63366[5:0] ^ p7_add_63366[10:5] ^ p7_add_63366[24:19], p7_add_63366[31:27] ^ p7_add_63366[4:0] ^ p7_add_63366[18:14], p7_add_63366[26:13] ^ p7_add_63366[31:18] ^ p7_add_63366[13:0], p7_add_63366[12:6] ^ p7_add_63366[17:11] ^ p7_add_63366[31:25]} + (p7_add_63366 & p7_add_63288 ^ ~(p7_add_63366 | ~p7_add_63212));
  assign p8_add_63447_comb = p7_message[255:227] + 29'h1b00_f553;
  assign p8_add_63443_comb = p8_add_63442_comb + p7_add_63370;
  assign p8_add_63470_comb = (p8_and_63451_comb ^ p7_add_63392 & p7_add_63238 ^ p7_and_63371) + p7_add_63365;
  assign p8_add_63444_comb = p8_add_63443_comb + p7_add_63238;
  assign p8_add_63450_comb = {p8_add_63447_comb, p7_message[226:224]} + p7_add_63212;
  assign p8_add_63472_comb = p8_add_63470_comb + {p7_add_63392[1:0] ^ p7_add_63392[12:11] ^ p7_add_63392[21:20], p7_add_63392[31:21] ^ p7_add_63392[10:0] ^ p7_add_63392[19:9], p7_add_63392[20:12] ^ p7_add_63392[31:23] ^ p7_add_63392[8:0], p7_add_63392[11:2] ^ p7_add_63392[22:13] ^ p7_add_63392[31:22]};

  // Registers for pipe stage 8:
  reg [511:0] p8_message;
  reg [31:0] p8_bit_slice_63040;
  reg [31:0] p8_bit_slice_63138;
  reg [31:0] p8_bit_slice_63213;
  reg [31:0] p8_add_63288;
  reg [31:0] p8_add_63366;
  reg [31:0] p8_bit_slice_63367;
  reg [31:0] p8_add_63443;
  reg [31:0] p8_add_63444;
  reg [31:0] p8_add_63450;
  reg [31:0] p8_add_63316;
  reg [31:0] p8_add_63392;
  reg [31:0] p8_and_63451;
  reg [31:0] p8_add_63472;
  always_ff @ (posedge clk) begin
    p8_message <= p7_message;
    p8_bit_slice_63040 <= p7_bit_slice_63040;
    p8_bit_slice_63138 <= p7_bit_slice_63138;
    p8_bit_slice_63213 <= p7_bit_slice_63213;
    p8_add_63288 <= p7_add_63288;
    p8_add_63366 <= p7_add_63366;
    p8_bit_slice_63367 <= p7_bit_slice_63367;
    p8_add_63443 <= p8_add_63443_comb;
    p8_add_63444 <= p8_add_63444_comb;
    p8_add_63450 <= p8_add_63450_comb;
    p8_add_63316 <= p7_add_63316;
    p8_add_63392 <= p7_add_63392;
    p8_and_63451 <= p8_and_63451_comb;
    p8_add_63472 <= p8_add_63472_comb;
  end

  // ===== Pipe stage 9:
  wire [31:0] p9_bit_slice_63525_comb;
  wire [31:0] p9_add_63584_comb;
  wire [31:0] p9_add_63585_comb;
  wire [31:0] p9_add_63586_comb;
  wire [31:0] p9_and_63529_comb;
  wire [31:0] p9_add_63522_comb;
  wire [31:0] p9_add_63523_comb;
  wire [31:0] p9_add_63527_comb;
  wire [31:0] p9_add_63548_comb;
  wire [31:0] p9_add_63524_comb;
  wire [31:0] p9_add_63528_comb;
  wire [31:0] p9_add_63550_comb;
  wire [31:0] p9_add_63603_comb;
  assign p9_bit_slice_63525_comb = p8_message[223:192];
  assign p9_add_63584_comb = p9_bit_slice_63525_comb + {p8_message[454:452] ^ p8_message[465:463], p8_message[451:448] ^ p8_message[462:459] ^ p8_message[479:476], p8_message[479:469] ^ p8_message[458:448] ^ p8_message[475:465], p8_message[468:455] ^ p8_message[479:466] ^ p8_message[464:451]};
  assign p9_add_63585_comb = {p8_message[48:39] ^ p8_message[50:41], p8_message[38:32] ^ p8_message[40:34] ^ p8_message[63:57], p8_message[63:62] ^ p8_message[33:32] ^ p8_message[56:55], p8_message[61:49] ^ p8_message[63:51] ^ p8_message[54:42]} + p8_message[511:480];
  assign p9_add_63586_comb = p9_add_63584_comb + p9_add_63585_comb;
  assign p9_and_63529_comb = p8_add_63472 & p8_add_63392;
  assign p9_add_63522_comb = (p8_add_63444 & p8_add_63366 ^ ~(p8_add_63444 | ~p8_add_63288)) + {p8_add_63444[5:0] ^ p8_add_63444[10:5] ^ p8_add_63444[24:19], p8_add_63444[31:27] ^ p8_add_63444[4:0] ^ p8_add_63444[18:14], p8_add_63444[26:13] ^ p8_add_63444[31:18] ^ p8_add_63444[13:0], p8_add_63444[12:6] ^ p8_add_63444[17:11] ^ p8_add_63444[31:25]};
  assign p9_add_63523_comb = p9_add_63522_comb + p8_add_63450;
  assign p9_add_63527_comb = p9_bit_slice_63525_comb + 32'h1283_5b01;
  assign p9_add_63548_comb = (p9_and_63529_comb ^ p8_add_63472 & p8_add_63316 ^ p8_and_63451) + p8_add_63443;
  assign p9_add_63524_comb = p9_add_63523_comb + p8_add_63316;
  assign p9_add_63528_comb = p8_add_63288 + p9_add_63527_comb;
  assign p9_add_63550_comb = p9_add_63548_comb + {p8_add_63472[1:0] ^ p8_add_63472[12:11] ^ p8_add_63472[21:20], p8_add_63472[31:21] ^ p8_add_63472[10:0] ^ p8_add_63472[19:9], p8_add_63472[20:12] ^ p8_add_63472[31:23] ^ p8_add_63472[8:0], p8_add_63472[11:2] ^ p8_add_63472[22:13] ^ p8_add_63472[31:22]};
  assign p9_add_63603_comb = {p9_add_63586_comb[16:7] ^ p9_add_63586_comb[18:9], p9_add_63586_comb[6:0] ^ p9_add_63586_comb[8:2] ^ p9_add_63586_comb[31:25], p9_add_63586_comb[31:30] ^ p9_add_63586_comb[1:0] ^ p9_add_63586_comb[24:23], p9_add_63586_comb[29:17] ^ p9_add_63586_comb[31:19] ^ p9_add_63586_comb[22:10]} + p8_bit_slice_63040;

  // Registers for pipe stage 9:
  reg [511:0] p9_message;
  reg [31:0] p9_bit_slice_63138;
  reg [31:0] p9_bit_slice_63213;
  reg [31:0] p9_add_63366;
  reg [31:0] p9_bit_slice_63367;
  reg [31:0] p9_add_63444;
  reg [31:0] p9_add_63523;
  reg [31:0] p9_add_63524;
  reg [31:0] p9_bit_slice_63525;
  reg [31:0] p9_add_63528;
  reg [31:0] p9_add_63392;
  reg [31:0] p9_add_63472;
  reg [31:0] p9_and_63529;
  reg [31:0] p9_add_63550;
  reg [31:0] p9_add_63586;
  reg [31:0] p9_add_63603;
  always_ff @ (posedge clk) begin
    p9_message <= p8_message;
    p9_bit_slice_63138 <= p8_bit_slice_63138;
    p9_bit_slice_63213 <= p8_bit_slice_63213;
    p9_add_63366 <= p8_add_63366;
    p9_bit_slice_63367 <= p8_bit_slice_63367;
    p9_add_63444 <= p8_add_63444;
    p9_add_63523 <= p9_add_63523_comb;
    p9_add_63524 <= p9_add_63524_comb;
    p9_bit_slice_63525 <= p9_bit_slice_63525_comb;
    p9_add_63528 <= p9_add_63528_comb;
    p9_add_63392 <= p8_add_63392;
    p9_add_63472 <= p8_add_63472;
    p9_and_63529 <= p9_and_63529_comb;
    p9_add_63550 <= p9_add_63550_comb;
    p9_add_63586 <= p9_add_63586_comb;
    p9_add_63603 <= p9_add_63603_comb;
  end

  // ===== Pipe stage 10:
  wire [31:0] p10_bit_slice_63666_comb;
  wire [31:0] p10_add_63742_comb;
  wire [1:0] p10_bit_slice_63689_comb;
  wire [31:0] p10_add_63743_comb;
  wire [31:0] p10_and_63667_comb;
  wire [31:0] p10_add_63657_comb;
  wire [30:0] p10_add_63662_comb;
  wire [31:0] p10_bit_slice_63719_comb;
  wire [31:0] p10_add_63658_comb;
  wire [31:0] p10_add_63686_comb;
  wire [31:0] p10_add_63723_comb;
  wire [31:0] p10_add_63724_comb;
  wire [31:0] p10_bit_slice_63774_comb;
  wire [31:0] p10_add_63659_comb;
  wire [31:0] p10_add_63665_comb;
  wire [31:0] p10_add_63688_comb;
  wire [31:0] p10_add_63725_comb;
  wire [31:0] p10_add_63777_comb;
  wire [31:0] p10_add_63778_comb;
  assign p10_bit_slice_63666_comb = p9_message[159:128];
  assign p10_add_63742_comb = p10_bit_slice_63666_comb + {p9_message[390:388] ^ p9_message[401:399], p9_message[387:384] ^ p9_message[398:395] ^ p9_message[415:412], p9_message[415:405] ^ p9_message[394:384] ^ p9_message[411:401], p9_message[404:391] ^ p9_message[415:402] ^ p9_message[400:387]};
  assign p10_bit_slice_63689_comb = p9_message[1:0];
  assign p10_add_63743_comb = p10_add_63742_comb + p9_add_63603;
  assign p10_and_63667_comb = p9_add_63550 & p9_add_63472;
  assign p10_add_63657_comb = {p9_add_63524[5:0] ^ p9_add_63524[10:5] ^ p9_add_63524[24:19], p9_add_63524[31:27] ^ p9_add_63524[4:0] ^ p9_add_63524[18:14], p9_add_63524[26:13] ^ p9_add_63524[31:18] ^ p9_add_63524[13:0], p9_add_63524[12:6] ^ p9_add_63524[17:11] ^ p9_add_63524[31:25]} + (p9_add_63524 & p9_add_63444 ^ ~(p9_add_63524 | ~p9_add_63366));
  assign p10_add_63662_comb = p9_message[191:161] + 31'h1218_c2df;
  assign p10_bit_slice_63719_comb = p9_message[191:160];
  assign p10_add_63658_comb = p10_add_63657_comb + p9_add_63528;
  assign p10_add_63686_comb = (p10_and_63667_comb ^ p9_add_63550 & p9_add_63392 ^ p9_and_63529) + p9_add_63523;
  assign p10_add_63723_comb = p10_bit_slice_63719_comb + {p9_message[422:420] ^ p9_message[433:431], p9_message[419:416] ^ p9_message[430:427] ^ p9_message[447:444], p9_message[447:437] ^ p9_message[426:416] ^ p9_message[443:433], p9_message[436:423] ^ p9_message[447:434] ^ p9_message[432:419]};
  assign p10_add_63724_comb = {p9_message[16:7] ^ p9_message[18:9], p9_message[6:0] ^ p9_message[8:2] ^ p9_message[31:25], p9_message[31:30] ^ p10_bit_slice_63689_comb ^ p9_message[24:23], p9_message[29:17] ^ p9_message[31:19] ^ p9_message[22:10]} + p9_message[479:448];
  assign p10_bit_slice_63774_comb = p9_message[95:64];
  assign p10_add_63659_comb = p10_add_63658_comb + p9_add_63392;
  assign p10_add_63665_comb = {p10_add_63662_comb, p9_message[160]} + p9_add_63366;
  assign p10_add_63688_comb = p10_add_63686_comb + {p9_add_63550[1:0] ^ p9_add_63550[12:11] ^ p9_add_63550[21:20], p9_add_63550[31:21] ^ p9_add_63550[10:0] ^ p9_add_63550[19:9], p9_add_63550[20:12] ^ p9_add_63550[31:23] ^ p9_add_63550[8:0], p9_add_63550[11:2] ^ p9_add_63550[22:13] ^ p9_add_63550[31:22]};
  assign p10_add_63725_comb = p10_add_63723_comb + p10_add_63724_comb;
  assign p10_add_63777_comb = p10_bit_slice_63774_comb + {p9_message[326:324] ^ p9_message[337:335], p9_message[323:320] ^ p9_message[334:331] ^ p9_message[351:348], p9_message[351:341] ^ p9_message[330:320] ^ p9_message[347:337], p9_message[340:327] ^ p9_message[351:338] ^ p9_message[336:323]};
  assign p10_add_63778_comb = {p10_add_63743_comb[16:7] ^ p10_add_63743_comb[18:9], p10_add_63743_comb[6:0] ^ p10_add_63743_comb[8:2] ^ p10_add_63743_comb[31:25], p10_add_63743_comb[31:30] ^ p10_add_63743_comb[1:0] ^ p10_add_63743_comb[24:23], p10_add_63743_comb[29:17] ^ p10_add_63743_comb[31:19] ^ p10_add_63743_comb[22:10]} + p9_bit_slice_63138;

  // Registers for pipe stage 10:
  reg [511:0] p10_message;
  reg [31:0] p10_bit_slice_63213;
  reg [31:0] p10_bit_slice_63367;
  reg [31:0] p10_add_63444;
  reg [31:0] p10_add_63524;
  reg [31:0] p10_bit_slice_63525;
  reg [31:0] p10_add_63658;
  reg [31:0] p10_add_63659;
  reg [31:0] p10_add_63665;
  reg [31:0] p10_add_63472;
  reg [31:0] p10_bit_slice_63666;
  reg [31:0] p10_add_63550;
  reg [31:0] p10_and_63667;
  reg [31:0] p10_add_63688;
  reg [1:0] p10_bit_slice_63689;
  reg [31:0] p10_add_63586;
  reg [31:0] p10_bit_slice_63719;
  reg [31:0] p10_add_63725;
  reg [31:0] p10_add_63743;
  reg [31:0] p10_bit_slice_63774;
  reg [31:0] p10_add_63777;
  reg [31:0] p10_add_63778;
  always_ff @ (posedge clk) begin
    p10_message <= p9_message;
    p10_bit_slice_63213 <= p9_bit_slice_63213;
    p10_bit_slice_63367 <= p9_bit_slice_63367;
    p10_add_63444 <= p9_add_63444;
    p10_add_63524 <= p9_add_63524;
    p10_bit_slice_63525 <= p9_bit_slice_63525;
    p10_add_63658 <= p10_add_63658_comb;
    p10_add_63659 <= p10_add_63659_comb;
    p10_add_63665 <= p10_add_63665_comb;
    p10_add_63472 <= p9_add_63472;
    p10_bit_slice_63666 <= p10_bit_slice_63666_comb;
    p10_add_63550 <= p9_add_63550;
    p10_and_63667 <= p10_and_63667_comb;
    p10_add_63688 <= p10_add_63688_comb;
    p10_bit_slice_63689 <= p10_bit_slice_63689_comb;
    p10_add_63586 <= p9_add_63586;
    p10_bit_slice_63719 <= p10_bit_slice_63719_comb;
    p10_add_63725 <= p10_add_63725_comb;
    p10_add_63743 <= p10_add_63743_comb;
    p10_bit_slice_63774 <= p10_bit_slice_63774_comb;
    p10_add_63777 <= p10_add_63777_comb;
    p10_add_63778 <= p10_add_63778_comb;
  end

  // ===== Pipe stage 11:
  wire [31:0] p11_bit_slice_63921_comb;
  wire [31:0] p11_add_63925_comb;
  wire [31:0] p11_add_63926_comb;
  wire [31:0] p11_add_63929_comb;
  wire [31:0] p11_add_63927_comb;
  wire [31:0] p11_add_63844_comb;
  wire [31:0] p11_and_63862_comb;
  wire [1:0] p11_bit_slice_63928_comb;
  wire [31:0] p11_add_63845_comb;
  wire [29:0] p11_add_63854_comb;
  wire [30:0] p11_add_63860_comb;
  wire [31:0] p11_bit_slice_63993_comb;
  wire [31:0] p11_add_63846_comb;
  wire [31:0] p11_add_63850_comb;
  wire [31:0] p11_add_63883_comb;
  wire [29:0] p11_add_63889_comb;
  wire [31:0] p11_bit_slice_63886_comb;
  wire [31:0] p11_add_63997_comb;
  wire [31:0] p11_add_63998_comb;
  wire [31:0] p11_nor_63848_comb;
  wire [31:0] p11_add_63851_comb;
  wire [31:0] p11_add_63857_comb;
  wire [31:0] p11_add_63882_comb;
  wire [31:0] p11_add_63885_comb;
  wire [31:0] p11_concat_63890_comb;
  wire [31:0] p11_add_63961_comb;
  wire [31:0] p11_add_63962_comb;
  wire [31:0] p11_add_63999_comb;
  wire [31:0] p11_add_64016_comb;
  wire [31:0] p11_bit_slice_64033_comb;
  wire [31:0] p11_add_64034_comb;
  wire [31:0] p11_add_64051_comb;
  wire [31:0] p11_add_64068_comb;
  wire [31:0] p11_add_64085_comb;
  wire [31:0] p11_concat_64101_comb;
  wire [31:0] p11_concat_64117_comb;
  wire [31:0] p11_concat_64133_comb;
  assign p11_bit_slice_63921_comb = p10_message[127:96];
  assign p11_add_63925_comb = p11_bit_slice_63921_comb + {p10_message[358:356] ^ p10_message[369:367], p10_message[355:352] ^ p10_message[366:363] ^ p10_message[383:380], p10_message[383:373] ^ p10_message[362:352] ^ p10_message[379:369], p10_message[372:359] ^ p10_message[383:370] ^ p10_message[368:355]};
  assign p11_add_63926_comb = {p10_add_63725[16:7] ^ p10_add_63725[18:9], p10_add_63725[6:0] ^ p10_add_63725[8:2] ^ p10_add_63725[31:25], p10_add_63725[31:30] ^ p10_add_63725[1:0] ^ p10_add_63725[24:23], p10_add_63725[29:17] ^ p10_add_63725[31:19] ^ p10_add_63725[22:10]} + p10_message[415:384];
  assign p11_add_63929_comb = p10_add_63777 + p10_add_63778;
  assign p11_add_63927_comb = p11_add_63925_comb + p11_add_63926_comb;
  assign p11_add_63844_comb = (p10_add_63659 & p10_add_63524 ^ ~(p10_add_63659 | ~p10_add_63444)) + {p10_add_63659[5:0] ^ p10_add_63659[10:5] ^ p10_add_63659[24:19], p10_add_63659[31:27] ^ p10_add_63659[4:0] ^ p10_add_63659[18:14], p10_add_63659[26:13] ^ p10_add_63659[31:18] ^ p10_add_63659[13:0], p10_add_63659[12:6] ^ p10_add_63659[17:11] ^ p10_add_63659[31:25]};
  assign p11_and_63862_comb = p10_add_63688 & p10_add_63550;
  assign p11_bit_slice_63928_comb = p11_add_63927_comb[1:0];
  assign p11_add_63845_comb = p11_add_63844_comb + p10_add_63665;
  assign p11_add_63854_comb = p10_message[127:98] + 30'h1caf_975d;
  assign p11_add_63860_comb = p10_message[95:65] + 31'h406f_58ff;
  assign p11_bit_slice_63993_comb = p10_message[31:0];
  assign p11_add_63846_comb = p11_add_63845_comb + p10_add_63472;
  assign p11_add_63850_comb = p10_bit_slice_63666 + 32'h550c_7dc3;
  assign p11_add_63883_comb = (p11_and_63862_comb ^ p10_add_63688 & p10_add_63472 ^ p10_and_63667) + p10_add_63658;
  assign p11_add_63889_comb = p10_message[31:2] + 30'h3066_fc5d;
  assign p11_bit_slice_63886_comb = p10_message[63:32];
  assign p11_add_63997_comb = p11_bit_slice_63993_comb + {p10_message[262:260] ^ p10_message[273:271], p10_message[259:256] ^ p10_message[270:267] ^ p10_message[287:284], p10_message[287:277] ^ p10_message[266:256] ^ p10_message[283:273], p10_message[276:263] ^ p10_message[287:274] ^ p10_message[272:259]};
  assign p11_add_63998_comb = {p11_add_63929_comb[16:7] ^ p11_add_63929_comb[18:9], p11_add_63929_comb[6:0] ^ p11_add_63929_comb[8:2] ^ p11_add_63929_comb[31:25], p11_add_63929_comb[31:30] ^ p11_add_63929_comb[1:0] ^ p11_add_63929_comb[24:23], p11_add_63929_comb[29:17] ^ p11_add_63929_comb[31:19] ^ p11_add_63929_comb[22:10]} + p10_message[319:288];
  assign p11_nor_63848_comb = ~(p11_add_63846_comb | ~p10_add_63524);
  assign p11_add_63851_comb = p10_add_63444 + p11_add_63850_comb;
  assign p11_add_63857_comb = {p11_add_63854_comb, p10_message[97:96]} + p10_add_63524;
  assign p11_add_63882_comb = {p11_add_63860_comb, p10_message[64]} + p10_add_63659;
  assign p11_add_63885_comb = p11_add_63883_comb + {p10_add_63688[1:0] ^ p10_add_63688[12:11] ^ p10_add_63688[21:20], p10_add_63688[31:21] ^ p10_add_63688[10:0] ^ p10_add_63688[19:9], p10_add_63688[20:12] ^ p10_add_63688[31:23] ^ p10_add_63688[8:0], p10_add_63688[11:2] ^ p10_add_63688[22:13] ^ p10_add_63688[31:22]};
  assign p11_concat_63890_comb = {p11_add_63889_comb, p10_bit_slice_63689};
  assign p11_add_63961_comb = p11_bit_slice_63886_comb + {p10_message[294:292] ^ p10_message[305:303], p10_message[291:288] ^ p10_message[302:299] ^ p10_message[319:316], p10_message[319:309] ^ p10_message[298:288] ^ p10_message[315:305], p10_message[308:295] ^ p10_message[319:306] ^ p10_message[304:291]};
  assign p11_add_63962_comb = {p11_add_63927_comb[16:7] ^ p11_add_63927_comb[18:9], p11_add_63927_comb[6:0] ^ p11_add_63927_comb[8:2] ^ p11_add_63927_comb[31:25], p11_add_63927_comb[31:30] ^ p11_bit_slice_63928_comb ^ p11_add_63927_comb[24:23], p11_add_63927_comb[29:17] ^ p11_add_63927_comb[31:19] ^ p11_add_63927_comb[22:10]} + p10_bit_slice_63213;
  assign p11_add_63999_comb = p11_add_63997_comb + p11_add_63998_comb;
  assign p11_add_64016_comb = p10_add_63586 + {p10_message[230:228] ^ p10_message[241:239], p10_message[227:224] ^ p10_message[238:235] ^ p10_message[255:252], p10_message[255:245] ^ p10_message[234:224] ^ p10_message[251:241], p10_message[244:231] ^ p10_message[255:242] ^ p10_message[240:227]};
  assign p11_bit_slice_64033_comb = p10_message[255:224];
  assign p11_add_64034_comb = p10_add_63725 + {p10_message[198:196] ^ p10_message[209:207], p10_message[195:192] ^ p10_message[206:203] ^ p10_message[223:220], p10_message[223:213] ^ p10_message[202:192] ^ p10_message[219:209], p10_message[212:199] ^ p10_message[223:210] ^ p10_message[208:195]};
  assign p11_add_64051_comb = p10_add_63743 + {p10_message[166:164] ^ p10_message[177:175], p10_message[163:160] ^ p10_message[174:171] ^ p10_message[191:188], p10_message[191:181] ^ p10_message[170:160] ^ p10_message[187:177], p10_message[180:167] ^ p10_message[191:178] ^ p10_message[176:163]};
  assign p11_add_64068_comb = p11_add_63927_comb + {p10_message[134:132] ^ p10_message[145:143], p10_message[131:128] ^ p10_message[142:139] ^ p10_message[159:156], p10_message[159:149] ^ p10_message[138:128] ^ p10_message[155:145], p10_message[148:135] ^ p10_message[159:146] ^ p10_message[144:131]};
  assign p11_add_64085_comb = p11_add_63929_comb + {p10_message[102:100] ^ p10_message[113:111], p10_message[99:96] ^ p10_message[110:107] ^ p10_message[127:124], p10_message[127:117] ^ p10_message[106:96] ^ p10_message[123:113], p10_message[116:103] ^ p10_message[127:114] ^ p10_message[112:99]};
  assign p11_concat_64101_comb = {p10_message[70:68] ^ p10_message[81:79], p10_message[67:64] ^ p10_message[78:75] ^ p10_message[95:92], p10_message[95:85] ^ p10_message[74:64] ^ p10_message[91:81], p10_message[84:71] ^ p10_message[95:82] ^ p10_message[80:67]};
  assign p11_concat_64117_comb = {p10_message[38:36] ^ p10_message[49:47], p10_message[35:32] ^ p10_message[46:43] ^ p10_message[63:60], p10_message[63:53] ^ p10_message[42:32] ^ p10_message[59:49], p10_message[52:39] ^ p10_message[63:50] ^ p10_message[48:35]};
  assign p11_concat_64133_comb = {p10_message[6:4] ^ p10_message[17:15], p10_message[3:0] ^ p10_message[14:11] ^ p10_message[31:28], p10_message[31:21] ^ p10_message[10:0] ^ p10_message[27:17], p10_message[20:7] ^ p10_message[31:18] ^ p10_message[16:3]};

  // Registers for pipe stage 11:
  reg [31:0] p11_bit_slice_63367;
  reg [31:0] p11_bit_slice_63525;
  reg [31:0] p11_add_63659;
  reg [31:0] p11_add_63845;
  reg [31:0] p11_add_63846;
  reg [31:0] p11_nor_63848;
  reg [31:0] p11_bit_slice_63666;
  reg [31:0] p11_add_63851;
  reg [31:0] p11_add_63550;
  reg [31:0] p11_add_63857;
  reg [31:0] p11_add_63688;
  reg [31:0] p11_and_63862;
  reg [31:0] p11_add_63882;
  reg [31:0] p11_add_63885;
  reg [31:0] p11_bit_slice_63886;
  reg [31:0] p11_concat_63890;
  reg [31:0] p11_add_63586;
  reg [31:0] p11_bit_slice_63719;
  reg [31:0] p11_add_63725;
  reg [31:0] p11_add_63743;
  reg [31:0] p11_bit_slice_63921;
  reg [31:0] p11_add_63927;
  reg [1:0] p11_bit_slice_63928;
  reg [31:0] p11_bit_slice_63774;
  reg [31:0] p11_add_63929;
  reg [31:0] p11_add_63961;
  reg [31:0] p11_add_63962;
  reg [31:0] p11_bit_slice_63993;
  reg [31:0] p11_add_63999;
  reg [31:0] p11_add_64016;
  reg [31:0] p11_bit_slice_64033;
  reg [31:0] p11_add_64034;
  reg [31:0] p11_add_64051;
  reg [31:0] p11_add_64068;
  reg [31:0] p11_add_64085;
  reg [31:0] p11_concat_64101;
  reg [31:0] p11_concat_64117;
  reg [31:0] p11_concat_64133;
  always_ff @ (posedge clk) begin
    p11_bit_slice_63367 <= p10_bit_slice_63367;
    p11_bit_slice_63525 <= p10_bit_slice_63525;
    p11_add_63659 <= p10_add_63659;
    p11_add_63845 <= p11_add_63845_comb;
    p11_add_63846 <= p11_add_63846_comb;
    p11_nor_63848 <= p11_nor_63848_comb;
    p11_bit_slice_63666 <= p10_bit_slice_63666;
    p11_add_63851 <= p11_add_63851_comb;
    p11_add_63550 <= p10_add_63550;
    p11_add_63857 <= p11_add_63857_comb;
    p11_add_63688 <= p10_add_63688;
    p11_and_63862 <= p11_and_63862_comb;
    p11_add_63882 <= p11_add_63882_comb;
    p11_add_63885 <= p11_add_63885_comb;
    p11_bit_slice_63886 <= p11_bit_slice_63886_comb;
    p11_concat_63890 <= p11_concat_63890_comb;
    p11_add_63586 <= p10_add_63586;
    p11_bit_slice_63719 <= p10_bit_slice_63719;
    p11_add_63725 <= p10_add_63725;
    p11_add_63743 <= p10_add_63743;
    p11_bit_slice_63921 <= p11_bit_slice_63921_comb;
    p11_add_63927 <= p11_add_63927_comb;
    p11_bit_slice_63928 <= p11_bit_slice_63928_comb;
    p11_bit_slice_63774 <= p10_bit_slice_63774;
    p11_add_63929 <= p11_add_63929_comb;
    p11_add_63961 <= p11_add_63961_comb;
    p11_add_63962 <= p11_add_63962_comb;
    p11_bit_slice_63993 <= p11_bit_slice_63993_comb;
    p11_add_63999 <= p11_add_63999_comb;
    p11_add_64016 <= p11_add_64016_comb;
    p11_bit_slice_64033 <= p11_bit_slice_64033_comb;
    p11_add_64034 <= p11_add_64034_comb;
    p11_add_64051 <= p11_add_64051_comb;
    p11_add_64068 <= p11_add_64068_comb;
    p11_add_64085 <= p11_add_64085_comb;
    p11_concat_64101 <= p11_concat_64101_comb;
    p11_concat_64117 <= p11_concat_64117_comb;
    p11_concat_64133 <= p11_concat_64133_comb;
  end

  // ===== Pipe stage 12:
  wire [1:0] p12_bit_slice_64257_comb;
  wire [31:0] p12_add_64256_comb;
  wire [31:0] p12_add_64291_comb;
  wire [31:0] p12_add_64292_comb;
  wire [31:0] p12_add_64229_comb;
  wire [31:0] p12_and_64234_comb;
  wire [31:0] p12_add_64230_comb;
  wire [31:0] p12_add_64231_comb;
  wire [31:0] p12_add_64253_comb;
  wire [31:0] p12_add_64274_comb;
  wire [31:0] p12_nor_64233_comb;
  wire [31:0] p12_add_64255_comb;
  wire [31:0] p12_add_64275_comb;
  wire [31:0] p12_add_64309_comb;
  wire [31:0] p12_add_64310_comb;
  wire [31:0] p12_add_64311_comb;
  assign p12_bit_slice_64257_comb = p11_add_63999[1:0];
  assign p12_add_64256_comb = p11_add_63961 + p11_add_63962;
  assign p12_add_64291_comb = {p11_add_63999[16:7] ^ p11_add_63999[18:9], p11_add_63999[6:0] ^ p11_add_63999[8:2] ^ p11_add_63999[31:25], p11_add_63999[31:30] ^ p12_bit_slice_64257_comb ^ p11_add_63999[24:23], p11_add_63999[29:17] ^ p11_add_63999[31:19] ^ p11_add_63999[22:10]} + p11_bit_slice_64033;
  assign p12_add_64292_comb = p11_add_64034 + p12_add_64291_comb;
  assign p12_add_64229_comb = {p11_add_63846[5:0] ^ p11_add_63846[10:5] ^ p11_add_63846[24:19], p11_add_63846[31:27] ^ p11_add_63846[4:0] ^ p11_add_63846[18:14], p11_add_63846[26:13] ^ p11_add_63846[31:18] ^ p11_add_63846[13:0], p11_add_63846[12:6] ^ p11_add_63846[17:11] ^ p11_add_63846[31:25]} + (p11_add_63846 & p11_add_63659 ^ p11_nor_63848);
  assign p12_and_64234_comb = p11_add_63885 & p11_add_63688;
  assign p12_add_64230_comb = p12_add_64229_comb + p11_add_63851;
  assign p12_add_64231_comb = p12_add_64230_comb + p11_add_63550;
  assign p12_add_64253_comb = (p12_and_64234_comb ^ p11_add_63885 & p11_add_63550 ^ p11_and_63862) + p11_add_63845;
  assign p12_add_64274_comb = {p12_add_64256_comb[16:7] ^ p12_add_64256_comb[18:9], p12_add_64256_comb[6:0] ^ p12_add_64256_comb[8:2] ^ p12_add_64256_comb[31:25], p12_add_64256_comb[31:30] ^ p12_add_64256_comb[1:0] ^ p12_add_64256_comb[24:23], p12_add_64256_comb[29:17] ^ p12_add_64256_comb[31:19] ^ p12_add_64256_comb[22:10]} + p11_bit_slice_63367;
  assign p12_nor_64233_comb = ~(p12_add_64231_comb | ~p11_add_63659);
  assign p12_add_64255_comb = p12_add_64253_comb + {p11_add_63885[1:0] ^ p11_add_63885[12:11] ^ p11_add_63885[21:20], p11_add_63885[31:21] ^ p11_add_63885[10:0] ^ p11_add_63885[19:9], p11_add_63885[20:12] ^ p11_add_63885[31:23] ^ p11_add_63885[8:0], p11_add_63885[11:2] ^ p11_add_63885[22:13] ^ p11_add_63885[31:22]};
  assign p12_add_64275_comb = p11_add_64016 + p12_add_64274_comb;
  assign p12_add_64309_comb = {p12_add_64292_comb[16:7] ^ p12_add_64292_comb[18:9], p12_add_64292_comb[6:0] ^ p12_add_64292_comb[8:2] ^ p12_add_64292_comb[31:25], p12_add_64292_comb[31:30] ^ p12_add_64292_comb[1:0] ^ p12_add_64292_comb[24:23], p12_add_64292_comb[29:17] ^ p12_add_64292_comb[31:19] ^ p12_add_64292_comb[22:10]} + p11_bit_slice_63719;
  assign p12_add_64310_comb = p12_add_64256_comb + p11_concat_64101;
  assign p12_add_64311_comb = p11_add_63999 + p11_concat_64117;

  // Registers for pipe stage 12:
  reg [31:0] p12_bit_slice_63525;
  reg [31:0] p12_add_63846;
  reg [31:0] p12_bit_slice_63666;
  reg [31:0] p12_add_64230;
  reg [31:0] p12_add_64231;
  reg [31:0] p12_nor_64233;
  reg [31:0] p12_add_63857;
  reg [31:0] p12_add_63688;
  reg [31:0] p12_add_63882;
  reg [31:0] p12_add_63885;
  reg [31:0] p12_bit_slice_63886;
  reg [31:0] p12_and_64234;
  reg [31:0] p12_add_64255;
  reg [31:0] p12_concat_63890;
  reg [31:0] p12_add_63586;
  reg [31:0] p12_add_63725;
  reg [31:0] p12_add_63743;
  reg [31:0] p12_bit_slice_63921;
  reg [31:0] p12_add_63927;
  reg [1:0] p12_bit_slice_63928;
  reg [31:0] p12_bit_slice_63774;
  reg [31:0] p12_add_63929;
  reg [31:0] p12_add_64256;
  reg [31:0] p12_bit_slice_63993;
  reg [31:0] p12_add_63999;
  reg [1:0] p12_bit_slice_64257;
  reg [31:0] p12_add_64275;
  reg [31:0] p12_add_64292;
  reg [31:0] p12_add_64051;
  reg [31:0] p12_add_64068;
  reg [31:0] p12_add_64309;
  reg [31:0] p12_add_64085;
  reg [31:0] p12_add_64310;
  reg [31:0] p12_add_64311;
  reg [31:0] p12_concat_64133;
  always_ff @ (posedge clk) begin
    p12_bit_slice_63525 <= p11_bit_slice_63525;
    p12_add_63846 <= p11_add_63846;
    p12_bit_slice_63666 <= p11_bit_slice_63666;
    p12_add_64230 <= p12_add_64230_comb;
    p12_add_64231 <= p12_add_64231_comb;
    p12_nor_64233 <= p12_nor_64233_comb;
    p12_add_63857 <= p11_add_63857;
    p12_add_63688 <= p11_add_63688;
    p12_add_63882 <= p11_add_63882;
    p12_add_63885 <= p11_add_63885;
    p12_bit_slice_63886 <= p11_bit_slice_63886;
    p12_and_64234 <= p12_and_64234_comb;
    p12_add_64255 <= p12_add_64255_comb;
    p12_concat_63890 <= p11_concat_63890;
    p12_add_63586 <= p11_add_63586;
    p12_add_63725 <= p11_add_63725;
    p12_add_63743 <= p11_add_63743;
    p12_bit_slice_63921 <= p11_bit_slice_63921;
    p12_add_63927 <= p11_add_63927;
    p12_bit_slice_63928 <= p11_bit_slice_63928;
    p12_bit_slice_63774 <= p11_bit_slice_63774;
    p12_add_63929 <= p11_add_63929;
    p12_add_64256 <= p12_add_64256_comb;
    p12_bit_slice_63993 <= p11_bit_slice_63993;
    p12_add_63999 <= p11_add_63999;
    p12_bit_slice_64257 <= p12_bit_slice_64257_comb;
    p12_add_64275 <= p12_add_64275_comb;
    p12_add_64292 <= p12_add_64292_comb;
    p12_add_64051 <= p11_add_64051;
    p12_add_64068 <= p11_add_64068;
    p12_add_64309 <= p12_add_64309_comb;
    p12_add_64085 <= p11_add_64085;
    p12_add_64310 <= p12_add_64310_comb;
    p12_add_64311 <= p12_add_64311_comb;
    p12_concat_64133 <= p11_concat_64133;
  end

  // ===== Pipe stage 13:
  wire [31:0] p13_add_64443_comb;
  wire [31:0] p13_add_64445_comb;
  wire [31:0] p13_add_64444_comb;
  wire [31:0] p13_and_64404_comb;
  wire [31:0] p13_add_64401_comb;
  wire [31:0] p13_add_64402_comb;
  wire [31:0] p13_add_64424_comb;
  wire [31:0] p13_add_64479_comb;
  wire [31:0] p13_add_64403_comb;
  wire [31:0] p13_add_64423_comb;
  wire [31:0] p13_add_64426_comb;
  wire [31:0] p13_add_64462_comb;
  wire [31:0] p13_add_64480_comb;
  wire [31:0] p13_add_64481_comb;
  assign p13_add_64443_comb = {p12_add_64275[16:7] ^ p12_add_64275[18:9], p12_add_64275[6:0] ^ p12_add_64275[8:2] ^ p12_add_64275[31:25], p12_add_64275[31:30] ^ p12_add_64275[1:0] ^ p12_add_64275[24:23], p12_add_64275[29:17] ^ p12_add_64275[31:19] ^ p12_add_64275[22:10]} + p12_bit_slice_63525;
  assign p13_add_64445_comb = p12_add_64068 + p12_add_64309;
  assign p13_add_64444_comb = p12_add_64051 + p13_add_64443_comb;
  assign p13_and_64404_comb = p12_add_64255 & p12_add_63885;
  assign p13_add_64401_comb = (p12_add_64231 & p12_add_63846 ^ p12_nor_64233) + {p12_add_64231[5:0] ^ p12_add_64231[10:5] ^ p12_add_64231[24:19], p12_add_64231[31:27] ^ p12_add_64231[4:0] ^ p12_add_64231[18:14], p12_add_64231[26:13] ^ p12_add_64231[31:18] ^ p12_add_64231[13:0], p12_add_64231[12:6] ^ p12_add_64231[17:11] ^ p12_add_64231[31:25]};
  assign p13_add_64402_comb = p13_add_64401_comb + p12_add_63857;
  assign p13_add_64424_comb = (p13_and_64404_comb ^ p12_add_64255 & p12_add_63688 ^ p12_and_64234) + p12_add_64230;
  assign p13_add_64479_comb = {p13_add_64445_comb[16:7] ^ p13_add_64445_comb[18:9], p13_add_64445_comb[6:0] ^ p13_add_64445_comb[8:2] ^ p13_add_64445_comb[31:25], p13_add_64445_comb[31:30] ^ p13_add_64445_comb[1:0] ^ p13_add_64445_comb[24:23], p13_add_64445_comb[29:17] ^ p13_add_64445_comb[31:19] ^ p13_add_64445_comb[22:10]} + p12_bit_slice_63921;
  assign p13_add_64403_comb = p13_add_64402_comb + p12_add_63688;
  assign p13_add_64423_comb = p12_concat_63890 + p12_add_64231;
  assign p13_add_64426_comb = p13_add_64424_comb + {p12_add_64255[1:0] ^ p12_add_64255[12:11] ^ p12_add_64255[21:20], p12_add_64255[31:21] ^ p12_add_64255[10:0] ^ p12_add_64255[19:9], p12_add_64255[20:12] ^ p12_add_64255[31:23] ^ p12_add_64255[8:0], p12_add_64255[11:2] ^ p12_add_64255[22:13] ^ p12_add_64255[31:22]};
  assign p13_add_64462_comb = {p13_add_64444_comb[16:7] ^ p13_add_64444_comb[18:9], p13_add_64444_comb[6:0] ^ p13_add_64444_comb[8:2] ^ p13_add_64444_comb[31:25], p13_add_64444_comb[31:30] ^ p13_add_64444_comb[1:0] ^ p13_add_64444_comb[24:23], p13_add_64444_comb[29:17] ^ p13_add_64444_comb[31:19] ^ p13_add_64444_comb[22:10]} + p12_bit_slice_63666;
  assign p13_add_64480_comb = p12_add_64310 + p13_add_64479_comb;
  assign p13_add_64481_comb = p12_add_64275 + p12_concat_64133;

  // Registers for pipe stage 13:
  reg [31:0] p13_add_63846;
  reg [31:0] p13_add_64231;
  reg [31:0] p13_add_64402;
  reg [31:0] p13_add_64403;
  reg [31:0] p13_add_63882;
  reg [31:0] p13_add_63885;
  reg [31:0] p13_bit_slice_63886;
  reg [31:0] p13_add_64255;
  reg [31:0] p13_and_64404;
  reg [31:0] p13_add_64423;
  reg [31:0] p13_add_64426;
  reg [31:0] p13_add_63586;
  reg [31:0] p13_add_63725;
  reg [31:0] p13_add_63743;
  reg [31:0] p13_add_63927;
  reg [1:0] p13_bit_slice_63928;
  reg [31:0] p13_bit_slice_63774;
  reg [31:0] p13_add_63929;
  reg [31:0] p13_add_64256;
  reg [31:0] p13_bit_slice_63993;
  reg [31:0] p13_add_63999;
  reg [1:0] p13_bit_slice_64257;
  reg [31:0] p13_add_64275;
  reg [31:0] p13_add_64292;
  reg [31:0] p13_add_64444;
  reg [31:0] p13_add_64445;
  reg [31:0] p13_add_64085;
  reg [31:0] p13_add_64462;
  reg [31:0] p13_add_64480;
  reg [31:0] p13_add_64311;
  reg [31:0] p13_add_64481;
  always_ff @ (posedge clk) begin
    p13_add_63846 <= p12_add_63846;
    p13_add_64231 <= p12_add_64231;
    p13_add_64402 <= p13_add_64402_comb;
    p13_add_64403 <= p13_add_64403_comb;
    p13_add_63882 <= p12_add_63882;
    p13_add_63885 <= p12_add_63885;
    p13_bit_slice_63886 <= p12_bit_slice_63886;
    p13_add_64255 <= p12_add_64255;
    p13_and_64404 <= p13_and_64404_comb;
    p13_add_64423 <= p13_add_64423_comb;
    p13_add_64426 <= p13_add_64426_comb;
    p13_add_63586 <= p12_add_63586;
    p13_add_63725 <= p12_add_63725;
    p13_add_63743 <= p12_add_63743;
    p13_add_63927 <= p12_add_63927;
    p13_bit_slice_63928 <= p12_bit_slice_63928;
    p13_bit_slice_63774 <= p12_bit_slice_63774;
    p13_add_63929 <= p12_add_63929;
    p13_add_64256 <= p12_add_64256;
    p13_bit_slice_63993 <= p12_bit_slice_63993;
    p13_add_63999 <= p12_add_63999;
    p13_bit_slice_64257 <= p12_bit_slice_64257;
    p13_add_64275 <= p12_add_64275;
    p13_add_64292 <= p12_add_64292;
    p13_add_64444 <= p13_add_64444_comb;
    p13_add_64445 <= p13_add_64445_comb;
    p13_add_64085 <= p12_add_64085;
    p13_add_64462 <= p13_add_64462_comb;
    p13_add_64480 <= p13_add_64480_comb;
    p13_add_64311 <= p12_add_64311;
    p13_add_64481 <= p13_add_64481_comb;
  end

  // ===== Pipe stage 14:
  wire [31:0] p14_add_64595_comb;
  wire [31:0] p14_add_64565_comb;
  wire [31:0] p14_and_64573_comb;
  wire [31:0] p14_add_64566_comb;
  wire [31:0] p14_add_64567_comb;
  wire [31:0] p14_add_64571_comb;
  wire [31:0] p14_add_64592_comb;
  wire [31:0] p14_add_64612_comb;
  wire [31:0] p14_add_64630_comb;
  wire [31:0] p14_nor_64569_comb;
  wire [31:0] p14_add_64572_comb;
  wire [31:0] p14_add_64594_comb;
  wire [31:0] p14_add_64613_comb;
  wire [31:0] p14_add_64631_comb;
  assign p14_add_64595_comb = p13_add_64085 + p13_add_64462;
  assign p14_add_64565_comb = (p13_add_64403 & p13_add_64231 ^ ~(p13_add_64403 | ~p13_add_63846)) + {p13_add_64403[5:0] ^ p13_add_64403[10:5] ^ p13_add_64403[24:19], p13_add_64403[31:27] ^ p13_add_64403[4:0] ^ p13_add_64403[18:14], p13_add_64403[26:13] ^ p13_add_64403[31:18] ^ p13_add_64403[13:0], p13_add_64403[12:6] ^ p13_add_64403[17:11] ^ p13_add_64403[31:25]};
  assign p14_and_64573_comb = p13_add_64426 & p13_add_64255;
  assign p14_add_64566_comb = p14_add_64565_comb + p13_add_63882;
  assign p14_add_64567_comb = p14_add_64566_comb + p13_add_63885;
  assign p14_add_64571_comb = p13_bit_slice_63886 + 32'h9bdc_06a7;
  assign p14_add_64592_comb = (p14_and_64573_comb ^ p13_add_64426 & p13_add_63885 ^ p13_and_64404) + p13_add_64402;
  assign p14_add_64612_comb = {p14_add_64595_comb[16:7] ^ p14_add_64595_comb[18:9], p14_add_64595_comb[6:0] ^ p14_add_64595_comb[8:2] ^ p14_add_64595_comb[31:25], p14_add_64595_comb[31:30] ^ p14_add_64595_comb[1:0] ^ p14_add_64595_comb[24:23], p14_add_64595_comb[29:17] ^ p14_add_64595_comb[31:19] ^ p14_add_64595_comb[22:10]} + p13_bit_slice_63774;
  assign p14_add_64630_comb = {p13_add_64480[16:7] ^ p13_add_64480[18:9], p13_add_64480[6:0] ^ p13_add_64480[8:2] ^ p13_add_64480[31:25], p13_add_64480[31:30] ^ p13_add_64480[1:0] ^ p13_add_64480[24:23], p13_add_64480[29:17] ^ p13_add_64480[31:19] ^ p13_add_64480[22:10]} + p13_bit_slice_63886;
  assign p14_nor_64569_comb = ~(p14_add_64567_comb | ~p13_add_64231);
  assign p14_add_64572_comb = p13_add_63846 + p14_add_64571_comb;
  assign p14_add_64594_comb = p14_add_64592_comb + {p13_add_64426[1:0] ^ p13_add_64426[12:11] ^ p13_add_64426[21:20], p13_add_64426[31:21] ^ p13_add_64426[10:0] ^ p13_add_64426[19:9], p13_add_64426[20:12] ^ p13_add_64426[31:23] ^ p13_add_64426[8:0], p13_add_64426[11:2] ^ p13_add_64426[22:13] ^ p13_add_64426[31:22]};
  assign p14_add_64613_comb = p13_add_64311 + p14_add_64612_comb;
  assign p14_add_64631_comb = p13_add_64481 + p14_add_64630_comb;

  // Registers for pipe stage 14:
  reg [31:0] p14_add_64403;
  reg [31:0] p14_add_64566;
  reg [31:0] p14_add_64567;
  reg [31:0] p14_nor_64569;
  reg [31:0] p14_add_64572;
  reg [31:0] p14_add_64255;
  reg [31:0] p14_add_64423;
  reg [31:0] p14_add_64426;
  reg [31:0] p14_add_63586;
  reg [31:0] p14_and_64573;
  reg [31:0] p14_add_64594;
  reg [31:0] p14_add_63725;
  reg [31:0] p14_add_63743;
  reg [31:0] p14_add_63927;
  reg [1:0] p14_bit_slice_63928;
  reg [31:0] p14_add_63929;
  reg [31:0] p14_add_64256;
  reg [31:0] p14_bit_slice_63993;
  reg [31:0] p14_add_63999;
  reg [1:0] p14_bit_slice_64257;
  reg [31:0] p14_add_64275;
  reg [31:0] p14_add_64292;
  reg [31:0] p14_add_64444;
  reg [31:0] p14_add_64445;
  reg [31:0] p14_add_64595;
  reg [31:0] p14_add_64480;
  reg [31:0] p14_add_64613;
  reg [31:0] p14_add_64631;
  always_ff @ (posedge clk) begin
    p14_add_64403 <= p13_add_64403;
    p14_add_64566 <= p14_add_64566_comb;
    p14_add_64567 <= p14_add_64567_comb;
    p14_nor_64569 <= p14_nor_64569_comb;
    p14_add_64572 <= p14_add_64572_comb;
    p14_add_64255 <= p13_add_64255;
    p14_add_64423 <= p13_add_64423;
    p14_add_64426 <= p13_add_64426;
    p14_add_63586 <= p13_add_63586;
    p14_and_64573 <= p14_and_64573_comb;
    p14_add_64594 <= p14_add_64594_comb;
    p14_add_63725 <= p13_add_63725;
    p14_add_63743 <= p13_add_63743;
    p14_add_63927 <= p13_add_63927;
    p14_bit_slice_63928 <= p13_bit_slice_63928;
    p14_add_63929 <= p13_add_63929;
    p14_add_64256 <= p13_add_64256;
    p14_bit_slice_63993 <= p13_bit_slice_63993;
    p14_add_63999 <= p13_add_63999;
    p14_bit_slice_64257 <= p13_bit_slice_64257;
    p14_add_64275 <= p13_add_64275;
    p14_add_64292 <= p13_add_64292;
    p14_add_64444 <= p13_add_64444;
    p14_add_64445 <= p13_add_64445;
    p14_add_64595 <= p14_add_64595_comb;
    p14_add_64480 <= p13_add_64480;
    p14_add_64613 <= p14_add_64613_comb;
    p14_add_64631 <= p14_add_64631_comb;
  end

  // ===== Pipe stage 15:
  wire [31:0] p15_and_64710_comb;
  wire [31:0] p15_add_64707_comb;
  wire [31:0] p15_add_64708_comb;
  wire [31:0] p15_add_64729_comb;
  wire [31:0] p15_add_64764_comb;
  wire [31:0] p15_add_64765_comb;
  wire [31:0] p15_add_64709_comb;
  wire [31:0] p15_add_64731_comb;
  wire [31:0] p15_add_64766_comb;
  assign p15_and_64710_comb = p14_add_64594 & p14_add_64426;
  assign p15_add_64707_comb = {p14_add_64567[5:0] ^ p14_add_64567[10:5] ^ p14_add_64567[24:19], p14_add_64567[31:27] ^ p14_add_64567[4:0] ^ p14_add_64567[18:14], p14_add_64567[26:13] ^ p14_add_64567[31:18] ^ p14_add_64567[13:0], p14_add_64567[12:6] ^ p14_add_64567[17:11] ^ p14_add_64567[31:25]} + (p14_add_64567 & p14_add_64403 ^ p14_nor_64569);
  assign p15_add_64708_comb = p15_add_64707_comb + p14_add_64572;
  assign p15_add_64729_comb = (p15_and_64710_comb ^ p14_add_64594 & p14_add_64255 ^ p14_and_64573) + p14_add_64566;
  assign p15_add_64764_comb = p14_add_64292 + {p14_add_63586[6:4] ^ p14_add_63586[17:15], p14_add_63586[3:0] ^ p14_add_63586[14:11] ^ p14_add_63586[31:28], p14_add_63586[31:21] ^ p14_add_63586[10:0] ^ p14_add_63586[27:17], p14_add_63586[20:7] ^ p14_add_63586[31:18] ^ p14_add_63586[16:3]};
  assign p15_add_64765_comb = {p14_add_64613[16:7] ^ p14_add_64613[18:9], p14_add_64613[6:0] ^ p14_add_64613[8:2] ^ p14_add_64613[31:25], p14_add_64613[31:30] ^ p14_add_64613[1:0] ^ p14_add_64613[24:23], p14_add_64613[29:17] ^ p14_add_64613[31:19] ^ p14_add_64613[22:10]} + p14_bit_slice_63993;
  assign p15_add_64709_comb = p15_add_64708_comb + p14_add_64255;
  assign p15_add_64731_comb = p15_add_64729_comb + {p14_add_64594[1:0] ^ p14_add_64594[12:11] ^ p14_add_64594[21:20], p14_add_64594[31:21] ^ p14_add_64594[10:0] ^ p14_add_64594[19:9], p14_add_64594[20:12] ^ p14_add_64594[31:23] ^ p14_add_64594[8:0], p14_add_64594[11:2] ^ p14_add_64594[22:13] ^ p14_add_64594[31:22]};
  assign p15_add_64766_comb = p15_add_64764_comb + p15_add_64765_comb;

  // Registers for pipe stage 15:
  reg [31:0] p15_add_64403;
  reg [31:0] p15_add_64567;
  reg [31:0] p15_add_64708;
  reg [31:0] p15_add_64709;
  reg [31:0] p15_add_64423;
  reg [31:0] p15_add_64426;
  reg [31:0] p15_add_63586;
  reg [31:0] p15_add_64594;
  reg [31:0] p15_add_63725;
  reg [31:0] p15_and_64710;
  reg [31:0] p15_add_64731;
  reg [31:0] p15_add_63743;
  reg [31:0] p15_add_63927;
  reg [1:0] p15_bit_slice_63928;
  reg [31:0] p15_add_63929;
  reg [31:0] p15_add_64256;
  reg [31:0] p15_add_63999;
  reg [1:0] p15_bit_slice_64257;
  reg [31:0] p15_add_64275;
  reg [31:0] p15_add_64292;
  reg [31:0] p15_add_64444;
  reg [31:0] p15_add_64445;
  reg [31:0] p15_add_64595;
  reg [31:0] p15_add_64480;
  reg [31:0] p15_add_64613;
  reg [31:0] p15_add_64631;
  reg [31:0] p15_add_64766;
  always_ff @ (posedge clk) begin
    p15_add_64403 <= p14_add_64403;
    p15_add_64567 <= p14_add_64567;
    p15_add_64708 <= p15_add_64708_comb;
    p15_add_64709 <= p15_add_64709_comb;
    p15_add_64423 <= p14_add_64423;
    p15_add_64426 <= p14_add_64426;
    p15_add_63586 <= p14_add_63586;
    p15_add_64594 <= p14_add_64594;
    p15_add_63725 <= p14_add_63725;
    p15_and_64710 <= p15_and_64710_comb;
    p15_add_64731 <= p15_add_64731_comb;
    p15_add_63743 <= p14_add_63743;
    p15_add_63927 <= p14_add_63927;
    p15_bit_slice_63928 <= p14_bit_slice_63928;
    p15_add_63929 <= p14_add_63929;
    p15_add_64256 <= p14_add_64256;
    p15_add_63999 <= p14_add_63999;
    p15_bit_slice_64257 <= p14_bit_slice_64257;
    p15_add_64275 <= p14_add_64275;
    p15_add_64292 <= p14_add_64292;
    p15_add_64444 <= p14_add_64444;
    p15_add_64445 <= p14_add_64445;
    p15_add_64595 <= p14_add_64595;
    p15_add_64480 <= p14_add_64480;
    p15_add_64613 <= p14_add_64613;
    p15_add_64631 <= p14_add_64631;
    p15_add_64766 <= p15_add_64766_comb;
  end

  // ===== Pipe stage 16:
  wire [31:0] p16_and_64848_comb;
  wire [31:0] p16_add_64842_comb;
  wire [31:0] p16_add_64843_comb;
  wire [31:0] p16_add_64846_comb;
  wire [31:0] p16_add_64867_comb;
  wire [31:0] p16_add_64902_comb;
  wire [31:0] p16_add_64903_comb;
  wire [31:0] p16_add_64844_comb;
  wire [31:0] p16_add_64847_comb;
  wire [31:0] p16_add_64869_comb;
  wire [31:0] p16_add_64904_comb;
  assign p16_and_64848_comb = p15_add_64731 & p15_add_64594;
  assign p16_add_64842_comb = (p15_add_64709 & p15_add_64567 ^ ~(p15_add_64709 | ~p15_add_64403)) + {p15_add_64709[5:0] ^ p15_add_64709[10:5] ^ p15_add_64709[24:19], p15_add_64709[31:27] ^ p15_add_64709[4:0] ^ p15_add_64709[18:14], p15_add_64709[26:13] ^ p15_add_64709[31:18] ^ p15_add_64709[13:0], p15_add_64709[12:6] ^ p15_add_64709[17:11] ^ p15_add_64709[31:25]};
  assign p16_add_64843_comb = p16_add_64842_comb + p15_add_64423;
  assign p16_add_64846_comb = p15_add_63586 + 32'he49b_69c1;
  assign p16_add_64867_comb = (p16_and_64848_comb ^ p15_add_64731 & p15_add_64426 ^ p15_and_64710) + p15_add_64708;
  assign p16_add_64902_comb = p15_add_64444 + {p15_add_63725[6:4] ^ p15_add_63725[17:15], p15_add_63725[3:0] ^ p15_add_63725[14:11] ^ p15_add_63725[31:28], p15_add_63725[31:21] ^ p15_add_63725[10:0] ^ p15_add_63725[27:17], p15_add_63725[20:7] ^ p15_add_63725[31:18] ^ p15_add_63725[16:3]};
  assign p16_add_64903_comb = {p15_add_64631[16:7] ^ p15_add_64631[18:9], p15_add_64631[6:0] ^ p15_add_64631[8:2] ^ p15_add_64631[31:25], p15_add_64631[31:30] ^ p15_add_64631[1:0] ^ p15_add_64631[24:23], p15_add_64631[29:17] ^ p15_add_64631[31:19] ^ p15_add_64631[22:10]} + p15_add_63586;
  assign p16_add_64844_comb = p16_add_64843_comb + p15_add_64426;
  assign p16_add_64847_comb = p15_add_64403 + p16_add_64846_comb;
  assign p16_add_64869_comb = p16_add_64867_comb + {p15_add_64731[1:0] ^ p15_add_64731[12:11] ^ p15_add_64731[21:20], p15_add_64731[31:21] ^ p15_add_64731[10:0] ^ p15_add_64731[19:9], p15_add_64731[20:12] ^ p15_add_64731[31:23] ^ p15_add_64731[8:0], p15_add_64731[11:2] ^ p15_add_64731[22:13] ^ p15_add_64731[31:22]};
  assign p16_add_64904_comb = p16_add_64902_comb + p16_add_64903_comb;

  // Registers for pipe stage 16:
  reg [31:0] p16_add_64567;
  reg [31:0] p16_add_64709;
  reg [31:0] p16_add_64843;
  reg [31:0] p16_add_64844;
  reg [31:0] p16_add_64847;
  reg [31:0] p16_add_64594;
  reg [31:0] p16_add_63725;
  reg [31:0] p16_add_64731;
  reg [31:0] p16_add_63743;
  reg [31:0] p16_and_64848;
  reg [31:0] p16_add_64869;
  reg [31:0] p16_add_63927;
  reg [1:0] p16_bit_slice_63928;
  reg [31:0] p16_add_63929;
  reg [31:0] p16_add_64256;
  reg [31:0] p16_add_63999;
  reg [1:0] p16_bit_slice_64257;
  reg [31:0] p16_add_64275;
  reg [31:0] p16_add_64292;
  reg [31:0] p16_add_64444;
  reg [31:0] p16_add_64445;
  reg [31:0] p16_add_64595;
  reg [31:0] p16_add_64480;
  reg [31:0] p16_add_64613;
  reg [31:0] p16_add_64631;
  reg [31:0] p16_add_64766;
  reg [31:0] p16_add_64904;
  always_ff @ (posedge clk) begin
    p16_add_64567 <= p15_add_64567;
    p16_add_64709 <= p15_add_64709;
    p16_add_64843 <= p16_add_64843_comb;
    p16_add_64844 <= p16_add_64844_comb;
    p16_add_64847 <= p16_add_64847_comb;
    p16_add_64594 <= p15_add_64594;
    p16_add_63725 <= p15_add_63725;
    p16_add_64731 <= p15_add_64731;
    p16_add_63743 <= p15_add_63743;
    p16_and_64848 <= p16_and_64848_comb;
    p16_add_64869 <= p16_add_64869_comb;
    p16_add_63927 <= p15_add_63927;
    p16_bit_slice_63928 <= p15_bit_slice_63928;
    p16_add_63929 <= p15_add_63929;
    p16_add_64256 <= p15_add_64256;
    p16_add_63999 <= p15_add_63999;
    p16_bit_slice_64257 <= p15_bit_slice_64257;
    p16_add_64275 <= p15_add_64275;
    p16_add_64292 <= p15_add_64292;
    p16_add_64444 <= p15_add_64444;
    p16_add_64445 <= p15_add_64445;
    p16_add_64595 <= p15_add_64595;
    p16_add_64480 <= p15_add_64480;
    p16_add_64613 <= p15_add_64613;
    p16_add_64631 <= p15_add_64631;
    p16_add_64766 <= p15_add_64766;
    p16_add_64904 <= p16_add_64904_comb;
  end

  // ===== Pipe stage 17:
  wire [31:0] p17_and_64989_comb;
  wire [31:0] p17_add_64980_comb;
  wire [30:0] p17_add_64985_comb;
  wire [31:0] p17_add_64981_comb;
  wire [31:0] p17_add_65008_comb;
  wire [31:0] p17_add_65043_comb;
  wire [31:0] p17_add_65044_comb;
  wire [31:0] p17_add_64982_comb;
  wire [31:0] p17_add_64988_comb;
  wire [31:0] p17_add_65010_comb;
  wire [31:0] p17_add_65045_comb;
  assign p17_and_64989_comb = p16_add_64869 & p16_add_64731;
  assign p17_add_64980_comb = {p16_add_64844[5:0] ^ p16_add_64844[10:5] ^ p16_add_64844[24:19], p16_add_64844[31:27] ^ p16_add_64844[4:0] ^ p16_add_64844[18:14], p16_add_64844[26:13] ^ p16_add_64844[31:18] ^ p16_add_64844[13:0], p16_add_64844[12:6] ^ p16_add_64844[17:11] ^ p16_add_64844[31:25]} + (p16_add_64844 & p16_add_64709 ^ ~(p16_add_64844 | ~p16_add_64567));
  assign p17_add_64985_comb = p16_add_63725[31:1] + 31'h77df_23c3;
  assign p17_add_64981_comb = p17_add_64980_comb + p16_add_64847;
  assign p17_add_65008_comb = (p17_and_64989_comb ^ p16_add_64869 & p16_add_64594 ^ p16_and_64848) + p16_add_64843;
  assign p17_add_65043_comb = p16_add_64445 + {p16_add_63743[6:4] ^ p16_add_63743[17:15], p16_add_63743[3:0] ^ p16_add_63743[14:11] ^ p16_add_63743[31:28], p16_add_63743[31:21] ^ p16_add_63743[10:0] ^ p16_add_63743[27:17], p16_add_63743[20:7] ^ p16_add_63743[31:18] ^ p16_add_63743[16:3]};
  assign p17_add_65044_comb = {p16_add_64766[16:7] ^ p16_add_64766[18:9], p16_add_64766[6:0] ^ p16_add_64766[8:2] ^ p16_add_64766[31:25], p16_add_64766[31:30] ^ p16_add_64766[1:0] ^ p16_add_64766[24:23], p16_add_64766[29:17] ^ p16_add_64766[31:19] ^ p16_add_64766[22:10]} + p16_add_63725;
  assign p17_add_64982_comb = p17_add_64981_comb + p16_add_64594;
  assign p17_add_64988_comb = {p17_add_64985_comb, p16_add_63725[0]} + p16_add_64567;
  assign p17_add_65010_comb = p17_add_65008_comb + {p16_add_64869[1:0] ^ p16_add_64869[12:11] ^ p16_add_64869[21:20], p16_add_64869[31:21] ^ p16_add_64869[10:0] ^ p16_add_64869[19:9], p16_add_64869[20:12] ^ p16_add_64869[31:23] ^ p16_add_64869[8:0], p16_add_64869[11:2] ^ p16_add_64869[22:13] ^ p16_add_64869[31:22]};
  assign p17_add_65045_comb = p17_add_65043_comb + p17_add_65044_comb;

  // Registers for pipe stage 17:
  reg [31:0] p17_add_64709;
  reg [31:0] p17_add_64844;
  reg [31:0] p17_add_64981;
  reg [31:0] p17_add_64982;
  reg [31:0] p17_add_64988;
  reg [31:0] p17_add_64731;
  reg [31:0] p17_add_63743;
  reg [31:0] p17_add_64869;
  reg [31:0] p17_add_63927;
  reg [1:0] p17_bit_slice_63928;
  reg [31:0] p17_and_64989;
  reg [31:0] p17_add_65010;
  reg [31:0] p17_add_63929;
  reg [31:0] p17_add_64256;
  reg [31:0] p17_add_63999;
  reg [1:0] p17_bit_slice_64257;
  reg [31:0] p17_add_64275;
  reg [31:0] p17_add_64292;
  reg [31:0] p17_add_64444;
  reg [31:0] p17_add_64445;
  reg [31:0] p17_add_64595;
  reg [31:0] p17_add_64480;
  reg [31:0] p17_add_64613;
  reg [31:0] p17_add_64631;
  reg [31:0] p17_add_64766;
  reg [31:0] p17_add_64904;
  reg [31:0] p17_add_65045;
  always_ff @ (posedge clk) begin
    p17_add_64709 <= p16_add_64709;
    p17_add_64844 <= p16_add_64844;
    p17_add_64981 <= p17_add_64981_comb;
    p17_add_64982 <= p17_add_64982_comb;
    p17_add_64988 <= p17_add_64988_comb;
    p17_add_64731 <= p16_add_64731;
    p17_add_63743 <= p16_add_63743;
    p17_add_64869 <= p16_add_64869;
    p17_add_63927 <= p16_add_63927;
    p17_bit_slice_63928 <= p16_bit_slice_63928;
    p17_and_64989 <= p17_and_64989_comb;
    p17_add_65010 <= p17_add_65010_comb;
    p17_add_63929 <= p16_add_63929;
    p17_add_64256 <= p16_add_64256;
    p17_add_63999 <= p16_add_63999;
    p17_bit_slice_64257 <= p16_bit_slice_64257;
    p17_add_64275 <= p16_add_64275;
    p17_add_64292 <= p16_add_64292;
    p17_add_64444 <= p16_add_64444;
    p17_add_64445 <= p16_add_64445;
    p17_add_64595 <= p16_add_64595;
    p17_add_64480 <= p16_add_64480;
    p17_add_64613 <= p16_add_64613;
    p17_add_64631 <= p16_add_64631;
    p17_add_64766 <= p16_add_64766;
    p17_add_64904 <= p16_add_64904;
    p17_add_65045 <= p17_add_65045_comb;
  end

  // ===== Pipe stage 18:
  wire [31:0] p18_and_65130_comb;
  wire [31:0] p18_add_65121_comb;
  wire [30:0] p18_add_65126_comb;
  wire [31:0] p18_add_65122_comb;
  wire [31:0] p18_add_65149_comb;
  wire [31:0] p18_add_65184_comb;
  wire [31:0] p18_add_65185_comb;
  wire [31:0] p18_add_65123_comb;
  wire [31:0] p18_add_65129_comb;
  wire [31:0] p18_add_65151_comb;
  wire [31:0] p18_add_65186_comb;
  assign p18_and_65130_comb = p17_add_65010 & p17_add_64869;
  assign p18_add_65121_comb = (p17_add_64982 & p17_add_64844 ^ ~(p17_add_64982 | ~p17_add_64709)) + {p17_add_64982[5:0] ^ p17_add_64982[10:5] ^ p17_add_64982[24:19], p17_add_64982[31:27] ^ p17_add_64982[4:0] ^ p17_add_64982[18:14], p17_add_64982[26:13] ^ p17_add_64982[31:18] ^ p17_add_64982[13:0], p17_add_64982[12:6] ^ p17_add_64982[17:11] ^ p17_add_64982[31:25]};
  assign p18_add_65126_comb = p17_add_63743[31:1] + 31'h07e0_cee3;
  assign p18_add_65122_comb = p18_add_65121_comb + p17_add_64988;
  assign p18_add_65149_comb = (p18_and_65130_comb ^ p17_add_65010 & p17_add_64731 ^ p17_and_64989) + p17_add_64981;
  assign p18_add_65184_comb = p17_add_64595 + {p17_add_63927[6:4] ^ p17_add_63927[17:15], p17_add_63927[3:0] ^ p17_add_63927[14:11] ^ p17_add_63927[31:28], p17_add_63927[31:21] ^ p17_add_63927[10:0] ^ p17_add_63927[27:17], p17_add_63927[20:7] ^ p17_add_63927[31:18] ^ p17_add_63927[16:3]};
  assign p18_add_65185_comb = {p17_add_64904[16:7] ^ p17_add_64904[18:9], p17_add_64904[6:0] ^ p17_add_64904[8:2] ^ p17_add_64904[31:25], p17_add_64904[31:30] ^ p17_add_64904[1:0] ^ p17_add_64904[24:23], p17_add_64904[29:17] ^ p17_add_64904[31:19] ^ p17_add_64904[22:10]} + p17_add_63743;
  assign p18_add_65123_comb = p18_add_65122_comb + p17_add_64731;
  assign p18_add_65129_comb = {p18_add_65126_comb, p17_add_63743[0]} + p17_add_64709;
  assign p18_add_65151_comb = p18_add_65149_comb + {p17_add_65010[1:0] ^ p17_add_65010[12:11] ^ p17_add_65010[21:20], p17_add_65010[31:21] ^ p17_add_65010[10:0] ^ p17_add_65010[19:9], p17_add_65010[20:12] ^ p17_add_65010[31:23] ^ p17_add_65010[8:0], p17_add_65010[11:2] ^ p17_add_65010[22:13] ^ p17_add_65010[31:22]};
  assign p18_add_65186_comb = p18_add_65184_comb + p18_add_65185_comb;

  // Registers for pipe stage 18:
  reg [31:0] p18_add_64844;
  reg [31:0] p18_add_64982;
  reg [31:0] p18_add_65122;
  reg [31:0] p18_add_65123;
  reg [31:0] p18_add_65129;
  reg [31:0] p18_add_64869;
  reg [31:0] p18_add_63927;
  reg [1:0] p18_bit_slice_63928;
  reg [31:0] p18_add_65010;
  reg [31:0] p18_add_63929;
  reg [31:0] p18_and_65130;
  reg [31:0] p18_add_65151;
  reg [31:0] p18_add_64256;
  reg [31:0] p18_add_63999;
  reg [1:0] p18_bit_slice_64257;
  reg [31:0] p18_add_64275;
  reg [31:0] p18_add_64292;
  reg [31:0] p18_add_64444;
  reg [31:0] p18_add_64445;
  reg [31:0] p18_add_64595;
  reg [31:0] p18_add_64480;
  reg [31:0] p18_add_64613;
  reg [31:0] p18_add_64631;
  reg [31:0] p18_add_64766;
  reg [31:0] p18_add_64904;
  reg [31:0] p18_add_65045;
  reg [31:0] p18_add_65186;
  always_ff @ (posedge clk) begin
    p18_add_64844 <= p17_add_64844;
    p18_add_64982 <= p17_add_64982;
    p18_add_65122 <= p18_add_65122_comb;
    p18_add_65123 <= p18_add_65123_comb;
    p18_add_65129 <= p18_add_65129_comb;
    p18_add_64869 <= p17_add_64869;
    p18_add_63927 <= p17_add_63927;
    p18_bit_slice_63928 <= p17_bit_slice_63928;
    p18_add_65010 <= p17_add_65010;
    p18_add_63929 <= p17_add_63929;
    p18_and_65130 <= p18_and_65130_comb;
    p18_add_65151 <= p18_add_65151_comb;
    p18_add_64256 <= p17_add_64256;
    p18_add_63999 <= p17_add_63999;
    p18_bit_slice_64257 <= p17_bit_slice_64257;
    p18_add_64275 <= p17_add_64275;
    p18_add_64292 <= p17_add_64292;
    p18_add_64444 <= p17_add_64444;
    p18_add_64445 <= p17_add_64445;
    p18_add_64595 <= p17_add_64595;
    p18_add_64480 <= p17_add_64480;
    p18_add_64613 <= p17_add_64613;
    p18_add_64631 <= p17_add_64631;
    p18_add_64766 <= p17_add_64766;
    p18_add_64904 <= p17_add_64904;
    p18_add_65045 <= p17_add_65045;
    p18_add_65186 <= p18_add_65186_comb;
  end

  // ===== Pipe stage 19:
  wire [31:0] p19_and_65270_comb;
  wire [31:0] p19_add_65262_comb;
  wire [29:0] p19_add_65267_comb;
  wire [31:0] p19_add_65263_comb;
  wire [31:0] p19_add_65289_comb;
  wire [31:0] p19_add_65324_comb;
  wire [31:0] p19_add_65325_comb;
  wire [31:0] p19_add_65264_comb;
  wire [31:0] p19_add_65269_comb;
  wire [31:0] p19_add_65291_comb;
  wire [31:0] p19_add_65326_comb;
  assign p19_and_65270_comb = p18_add_65151 & p18_add_65010;
  assign p19_add_65262_comb = (p18_add_65123 & p18_add_64982 ^ ~(p18_add_65123 | ~p18_add_64844)) + {p18_add_65123[5:0] ^ p18_add_65123[10:5] ^ p18_add_65123[24:19], p18_add_65123[31:27] ^ p18_add_65123[4:0] ^ p18_add_65123[18:14], p18_add_65123[26:13] ^ p18_add_65123[31:18] ^ p18_add_65123[13:0], p18_add_65123[12:6] ^ p18_add_65123[17:11] ^ p18_add_65123[31:25]};
  assign p19_add_65267_comb = p18_add_63927[31:2] + 30'h0903_2873;
  assign p19_add_65263_comb = p19_add_65262_comb + p18_add_65129;
  assign p19_add_65289_comb = (p19_and_65270_comb ^ p18_add_65151 & p18_add_64869 ^ p18_and_65130) + p18_add_65122;
  assign p19_add_65324_comb = p18_add_64480 + {p18_add_63929[6:4] ^ p18_add_63929[17:15], p18_add_63929[3:0] ^ p18_add_63929[14:11] ^ p18_add_63929[31:28], p18_add_63929[31:21] ^ p18_add_63929[10:0] ^ p18_add_63929[27:17], p18_add_63929[20:7] ^ p18_add_63929[31:18] ^ p18_add_63929[16:3]};
  assign p19_add_65325_comb = {p18_add_65045[16:7] ^ p18_add_65045[18:9], p18_add_65045[6:0] ^ p18_add_65045[8:2] ^ p18_add_65045[31:25], p18_add_65045[31:30] ^ p18_add_65045[1:0] ^ p18_add_65045[24:23], p18_add_65045[29:17] ^ p18_add_65045[31:19] ^ p18_add_65045[22:10]} + p18_add_63927;
  assign p19_add_65264_comb = p19_add_65263_comb + p18_add_64869;
  assign p19_add_65269_comb = {p19_add_65267_comb, p18_bit_slice_63928} + p18_add_64844;
  assign p19_add_65291_comb = p19_add_65289_comb + {p18_add_65151[1:0] ^ p18_add_65151[12:11] ^ p18_add_65151[21:20], p18_add_65151[31:21] ^ p18_add_65151[10:0] ^ p18_add_65151[19:9], p18_add_65151[20:12] ^ p18_add_65151[31:23] ^ p18_add_65151[8:0], p18_add_65151[11:2] ^ p18_add_65151[22:13] ^ p18_add_65151[31:22]};
  assign p19_add_65326_comb = p19_add_65324_comb + p19_add_65325_comb;

  // Registers for pipe stage 19:
  reg [31:0] p19_add_64982;
  reg [31:0] p19_add_65123;
  reg [31:0] p19_add_65263;
  reg [31:0] p19_add_65264;
  reg [31:0] p19_add_65269;
  reg [31:0] p19_add_65010;
  reg [31:0] p19_add_63929;
  reg [31:0] p19_add_65151;
  reg [31:0] p19_add_64256;
  reg [31:0] p19_and_65270;
  reg [31:0] p19_add_65291;
  reg [31:0] p19_add_63999;
  reg [1:0] p19_bit_slice_64257;
  reg [31:0] p19_add_64275;
  reg [31:0] p19_add_64292;
  reg [31:0] p19_add_64444;
  reg [31:0] p19_add_64445;
  reg [31:0] p19_add_64595;
  reg [31:0] p19_add_64480;
  reg [31:0] p19_add_64613;
  reg [31:0] p19_add_64631;
  reg [31:0] p19_add_64766;
  reg [31:0] p19_add_64904;
  reg [31:0] p19_add_65045;
  reg [31:0] p19_add_65186;
  reg [31:0] p19_add_65326;
  always_ff @ (posedge clk) begin
    p19_add_64982 <= p18_add_64982;
    p19_add_65123 <= p18_add_65123;
    p19_add_65263 <= p19_add_65263_comb;
    p19_add_65264 <= p19_add_65264_comb;
    p19_add_65269 <= p19_add_65269_comb;
    p19_add_65010 <= p18_add_65010;
    p19_add_63929 <= p18_add_63929;
    p19_add_65151 <= p18_add_65151;
    p19_add_64256 <= p18_add_64256;
    p19_and_65270 <= p19_and_65270_comb;
    p19_add_65291 <= p19_add_65291_comb;
    p19_add_63999 <= p18_add_63999;
    p19_bit_slice_64257 <= p18_bit_slice_64257;
    p19_add_64275 <= p18_add_64275;
    p19_add_64292 <= p18_add_64292;
    p19_add_64444 <= p18_add_64444;
    p19_add_64445 <= p18_add_64445;
    p19_add_64595 <= p18_add_64595;
    p19_add_64480 <= p18_add_64480;
    p19_add_64613 <= p18_add_64613;
    p19_add_64631 <= p18_add_64631;
    p19_add_64766 <= p18_add_64766;
    p19_add_64904 <= p18_add_64904;
    p19_add_65045 <= p18_add_65045;
    p19_add_65186 <= p18_add_65186;
    p19_add_65326 <= p19_add_65326_comb;
  end

  // ===== Pipe stage 20:
  wire [31:0] p20_and_65406_comb;
  wire [31:0] p20_add_65400_comb;
  wire [31:0] p20_add_65401_comb;
  wire [31:0] p20_add_65404_comb;
  wire [31:0] p20_add_65425_comb;
  wire [31:0] p20_add_65402_comb;
  wire [31:0] p20_add_65405_comb;
  wire [31:0] p20_add_65427_comb;
  assign p20_and_65406_comb = p19_add_65291 & p19_add_65151;
  assign p20_add_65400_comb = (p19_add_65264 & p19_add_65123 ^ ~(p19_add_65264 | ~p19_add_64982)) + {p19_add_65264[5:0] ^ p19_add_65264[10:5] ^ p19_add_65264[24:19], p19_add_65264[31:27] ^ p19_add_65264[4:0] ^ p19_add_65264[18:14], p19_add_65264[26:13] ^ p19_add_65264[31:18] ^ p19_add_65264[13:0], p19_add_65264[12:6] ^ p19_add_65264[17:11] ^ p19_add_65264[31:25]};
  assign p20_add_65401_comb = p20_add_65400_comb + p19_add_65269;
  assign p20_add_65404_comb = p19_add_63929 + 32'h2de9_2c6f;
  assign p20_add_65425_comb = (p20_and_65406_comb ^ p19_add_65291 & p19_add_65010 ^ p19_and_65270) + p19_add_65263;
  assign p20_add_65402_comb = p20_add_65401_comb + p19_add_65010;
  assign p20_add_65405_comb = p19_add_64982 + p20_add_65404_comb;
  assign p20_add_65427_comb = p20_add_65425_comb + {p19_add_65291[1:0] ^ p19_add_65291[12:11] ^ p19_add_65291[21:20], p19_add_65291[31:21] ^ p19_add_65291[10:0] ^ p19_add_65291[19:9], p19_add_65291[20:12] ^ p19_add_65291[31:23] ^ p19_add_65291[8:0], p19_add_65291[11:2] ^ p19_add_65291[22:13] ^ p19_add_65291[31:22]};

  // Registers for pipe stage 20:
  reg [31:0] p20_add_65123;
  reg [31:0] p20_add_65264;
  reg [31:0] p20_add_65401;
  reg [31:0] p20_add_65402;
  reg [31:0] p20_add_63929;
  reg [31:0] p20_add_65405;
  reg [31:0] p20_add_65151;
  reg [31:0] p20_add_64256;
  reg [31:0] p20_add_65291;
  reg [31:0] p20_add_63999;
  reg [1:0] p20_bit_slice_64257;
  reg [31:0] p20_and_65406;
  reg [31:0] p20_add_65427;
  reg [31:0] p20_add_64275;
  reg [31:0] p20_add_64292;
  reg [31:0] p20_add_64444;
  reg [31:0] p20_add_64445;
  reg [31:0] p20_add_64595;
  reg [31:0] p20_add_64480;
  reg [31:0] p20_add_64613;
  reg [31:0] p20_add_64631;
  reg [31:0] p20_add_64766;
  reg [31:0] p20_add_64904;
  reg [31:0] p20_add_65045;
  reg [31:0] p20_add_65186;
  reg [31:0] p20_add_65326;
  always_ff @ (posedge clk) begin
    p20_add_65123 <= p19_add_65123;
    p20_add_65264 <= p19_add_65264;
    p20_add_65401 <= p20_add_65401_comb;
    p20_add_65402 <= p20_add_65402_comb;
    p20_add_63929 <= p19_add_63929;
    p20_add_65405 <= p20_add_65405_comb;
    p20_add_65151 <= p19_add_65151;
    p20_add_64256 <= p19_add_64256;
    p20_add_65291 <= p19_add_65291;
    p20_add_63999 <= p19_add_63999;
    p20_bit_slice_64257 <= p19_bit_slice_64257;
    p20_and_65406 <= p20_and_65406_comb;
    p20_add_65427 <= p20_add_65427_comb;
    p20_add_64275 <= p19_add_64275;
    p20_add_64292 <= p19_add_64292;
    p20_add_64444 <= p19_add_64444;
    p20_add_64445 <= p19_add_64445;
    p20_add_64595 <= p19_add_64595;
    p20_add_64480 <= p19_add_64480;
    p20_add_64613 <= p19_add_64613;
    p20_add_64631 <= p19_add_64631;
    p20_add_64766 <= p19_add_64766;
    p20_add_64904 <= p19_add_64904;
    p20_add_65045 <= p19_add_65045;
    p20_add_65186 <= p19_add_65186;
    p20_add_65326 <= p19_add_65326;
  end

  // ===== Pipe stage 21:
  wire [31:0] p21_and_65510_comb;
  wire [31:0] p21_add_65501_comb;
  wire [30:0] p21_add_65506_comb;
  wire [31:0] p21_add_65502_comb;
  wire [31:0] p21_add_65529_comb;
  wire [31:0] p21_add_65503_comb;
  wire [31:0] p21_add_65509_comb;
  wire [31:0] p21_add_65531_comb;
  assign p21_and_65510_comb = p20_add_65427 & p20_add_65291;
  assign p21_add_65501_comb = {p20_add_65402[5:0] ^ p20_add_65402[10:5] ^ p20_add_65402[24:19], p20_add_65402[31:27] ^ p20_add_65402[4:0] ^ p20_add_65402[18:14], p20_add_65402[26:13] ^ p20_add_65402[31:18] ^ p20_add_65402[13:0], p20_add_65402[12:6] ^ p20_add_65402[17:11] ^ p20_add_65402[31:25]} + (p20_add_65402 & p20_add_65264 ^ ~(p20_add_65402 | ~p20_add_65123));
  assign p21_add_65506_comb = p20_add_64256[31:1] + 31'h253a_4255;
  assign p21_add_65502_comb = p21_add_65501_comb + p20_add_65405;
  assign p21_add_65529_comb = (p21_and_65510_comb ^ p20_add_65427 & p20_add_65151 ^ p20_and_65406) + p20_add_65401;
  assign p21_add_65503_comb = p21_add_65502_comb + p20_add_65151;
  assign p21_add_65509_comb = {p21_add_65506_comb, p20_add_64256[0]} + p20_add_65123;
  assign p21_add_65531_comb = p21_add_65529_comb + {p20_add_65427[1:0] ^ p20_add_65427[12:11] ^ p20_add_65427[21:20], p20_add_65427[31:21] ^ p20_add_65427[10:0] ^ p20_add_65427[19:9], p20_add_65427[20:12] ^ p20_add_65427[31:23] ^ p20_add_65427[8:0], p20_add_65427[11:2] ^ p20_add_65427[22:13] ^ p20_add_65427[31:22]};

  // Registers for pipe stage 21:
  reg [31:0] p21_add_65264;
  reg [31:0] p21_add_65402;
  reg [31:0] p21_add_63929;
  reg [31:0] p21_add_65502;
  reg [31:0] p21_add_65503;
  reg [31:0] p21_add_64256;
  reg [31:0] p21_add_65509;
  reg [31:0] p21_add_65291;
  reg [31:0] p21_add_63999;
  reg [1:0] p21_bit_slice_64257;
  reg [31:0] p21_add_65427;
  reg [31:0] p21_add_64275;
  reg [31:0] p21_and_65510;
  reg [31:0] p21_add_65531;
  reg [31:0] p21_add_64292;
  reg [31:0] p21_add_64444;
  reg [31:0] p21_add_64445;
  reg [31:0] p21_add_64595;
  reg [31:0] p21_add_64480;
  reg [31:0] p21_add_64613;
  reg [31:0] p21_add_64631;
  reg [31:0] p21_add_64766;
  reg [31:0] p21_add_64904;
  reg [31:0] p21_add_65045;
  reg [31:0] p21_add_65186;
  reg [31:0] p21_add_65326;
  always_ff @ (posedge clk) begin
    p21_add_65264 <= p20_add_65264;
    p21_add_65402 <= p20_add_65402;
    p21_add_63929 <= p20_add_63929;
    p21_add_65502 <= p21_add_65502_comb;
    p21_add_65503 <= p21_add_65503_comb;
    p21_add_64256 <= p20_add_64256;
    p21_add_65509 <= p21_add_65509_comb;
    p21_add_65291 <= p20_add_65291;
    p21_add_63999 <= p20_add_63999;
    p21_bit_slice_64257 <= p20_bit_slice_64257;
    p21_add_65427 <= p20_add_65427;
    p21_add_64275 <= p20_add_64275;
    p21_and_65510 <= p21_and_65510_comb;
    p21_add_65531 <= p21_add_65531_comb;
    p21_add_64292 <= p20_add_64292;
    p21_add_64444 <= p20_add_64444;
    p21_add_64445 <= p20_add_64445;
    p21_add_64595 <= p20_add_64595;
    p21_add_64480 <= p20_add_64480;
    p21_add_64613 <= p20_add_64613;
    p21_add_64631 <= p20_add_64631;
    p21_add_64766 <= p20_add_64766;
    p21_add_64904 <= p20_add_64904;
    p21_add_65045 <= p20_add_65045;
    p21_add_65186 <= p20_add_65186;
    p21_add_65326 <= p20_add_65326;
  end

  // ===== Pipe stage 22:
  wire [31:0] p22_and_65613_comb;
  wire [31:0] p22_add_65605_comb;
  wire [29:0] p22_add_65610_comb;
  wire [31:0] p22_add_65606_comb;
  wire [31:0] p22_add_65632_comb;
  wire [31:0] p22_add_65607_comb;
  wire [31:0] p22_add_65612_comb;
  wire [31:0] p22_add_65634_comb;
  assign p22_and_65613_comb = p21_add_65531 & p21_add_65427;
  assign p22_add_65605_comb = (p21_add_65503 & p21_add_65402 ^ ~(p21_add_65503 | ~p21_add_65264)) + {p21_add_65503[5:0] ^ p21_add_65503[10:5] ^ p21_add_65503[24:19], p21_add_65503[31:27] ^ p21_add_65503[4:0] ^ p21_add_65503[18:14], p21_add_65503[26:13] ^ p21_add_65503[31:18] ^ p21_add_65503[13:0], p21_add_65503[12:6] ^ p21_add_65503[17:11] ^ p21_add_65503[31:25]};
  assign p22_add_65610_comb = p21_add_63999[31:2] + 30'h172c_2a77;
  assign p22_add_65606_comb = p22_add_65605_comb + p21_add_65509;
  assign p22_add_65632_comb = (p22_and_65613_comb ^ p21_add_65531 & p21_add_65291 ^ p21_and_65510) + p21_add_65502;
  assign p22_add_65607_comb = p22_add_65606_comb + p21_add_65291;
  assign p22_add_65612_comb = {p22_add_65610_comb, p21_bit_slice_64257} + p21_add_65264;
  assign p22_add_65634_comb = p22_add_65632_comb + {p21_add_65531[1:0] ^ p21_add_65531[12:11] ^ p21_add_65531[21:20], p21_add_65531[31:21] ^ p21_add_65531[10:0] ^ p21_add_65531[19:9], p21_add_65531[20:12] ^ p21_add_65531[31:23] ^ p21_add_65531[8:0], p21_add_65531[11:2] ^ p21_add_65531[22:13] ^ p21_add_65531[31:22]};

  // Registers for pipe stage 22:
  reg [31:0] p22_add_65402;
  reg [31:0] p22_add_63929;
  reg [31:0] p22_add_65503;
  reg [31:0] p22_add_64256;
  reg [31:0] p22_add_65606;
  reg [31:0] p22_add_65607;
  reg [31:0] p22_add_63999;
  reg [31:0] p22_add_65612;
  reg [31:0] p22_add_65427;
  reg [31:0] p22_add_64275;
  reg [31:0] p22_add_65531;
  reg [31:0] p22_add_64292;
  reg [31:0] p22_and_65613;
  reg [31:0] p22_add_65634;
  reg [31:0] p22_add_64444;
  reg [31:0] p22_add_64445;
  reg [31:0] p22_add_64595;
  reg [31:0] p22_add_64480;
  reg [31:0] p22_add_64613;
  reg [31:0] p22_add_64631;
  reg [31:0] p22_add_64766;
  reg [31:0] p22_add_64904;
  reg [31:0] p22_add_65045;
  reg [31:0] p22_add_65186;
  reg [31:0] p22_add_65326;
  always_ff @ (posedge clk) begin
    p22_add_65402 <= p21_add_65402;
    p22_add_63929 <= p21_add_63929;
    p22_add_65503 <= p21_add_65503;
    p22_add_64256 <= p21_add_64256;
    p22_add_65606 <= p22_add_65606_comb;
    p22_add_65607 <= p22_add_65607_comb;
    p22_add_63999 <= p21_add_63999;
    p22_add_65612 <= p22_add_65612_comb;
    p22_add_65427 <= p21_add_65427;
    p22_add_64275 <= p21_add_64275;
    p22_add_65531 <= p21_add_65531;
    p22_add_64292 <= p21_add_64292;
    p22_and_65613 <= p22_and_65613_comb;
    p22_add_65634 <= p22_add_65634_comb;
    p22_add_64444 <= p21_add_64444;
    p22_add_64445 <= p21_add_64445;
    p22_add_64595 <= p21_add_64595;
    p22_add_64480 <= p21_add_64480;
    p22_add_64613 <= p21_add_64613;
    p22_add_64631 <= p21_add_64631;
    p22_add_64766 <= p21_add_64766;
    p22_add_64904 <= p21_add_64904;
    p22_add_65045 <= p21_add_65045;
    p22_add_65186 <= p21_add_65186;
    p22_add_65326 <= p21_add_65326;
  end

  // ===== Pipe stage 23:
  wire [31:0] p23_and_65715_comb;
  wire [31:0] p23_add_65706_comb;
  wire [30:0] p23_add_65711_comb;
  wire [31:0] p23_add_65707_comb;
  wire [31:0] p23_add_65734_comb;
  wire [31:0] p23_add_65708_comb;
  wire [31:0] p23_add_65714_comb;
  wire [31:0] p23_add_65736_comb;
  assign p23_and_65715_comb = p22_add_65634 & p22_add_65531;
  assign p23_add_65706_comb = (p22_add_65607 & p22_add_65503 ^ ~(p22_add_65607 | ~p22_add_65402)) + {p22_add_65607[5:0] ^ p22_add_65607[10:5] ^ p22_add_65607[24:19], p22_add_65607[31:27] ^ p22_add_65607[4:0] ^ p22_add_65607[18:14], p22_add_65607[26:13] ^ p22_add_65607[31:18] ^ p22_add_65607[13:0], p22_add_65607[12:6] ^ p22_add_65607[17:11] ^ p22_add_65607[31:25]};
  assign p23_add_65711_comb = p22_add_64275[31:1] + 31'h3b7c_c46d;
  assign p23_add_65707_comb = p23_add_65706_comb + p22_add_65612;
  assign p23_add_65734_comb = (p23_and_65715_comb ^ p22_add_65634 & p22_add_65427 ^ p22_and_65613) + p22_add_65606;
  assign p23_add_65708_comb = p23_add_65707_comb + p22_add_65427;
  assign p23_add_65714_comb = {p23_add_65711_comb, p22_add_64275[0]} + p22_add_65402;
  assign p23_add_65736_comb = p23_add_65734_comb + {p22_add_65634[1:0] ^ p22_add_65634[12:11] ^ p22_add_65634[21:20], p22_add_65634[31:21] ^ p22_add_65634[10:0] ^ p22_add_65634[19:9], p22_add_65634[20:12] ^ p22_add_65634[31:23] ^ p22_add_65634[8:0], p22_add_65634[11:2] ^ p22_add_65634[22:13] ^ p22_add_65634[31:22]};

  // Registers for pipe stage 23:
  reg [31:0] p23_add_63929;
  reg [31:0] p23_add_65503;
  reg [31:0] p23_add_64256;
  reg [31:0] p23_add_65607;
  reg [31:0] p23_add_63999;
  reg [31:0] p23_add_65707;
  reg [31:0] p23_add_65708;
  reg [31:0] p23_add_64275;
  reg [31:0] p23_add_65714;
  reg [31:0] p23_add_65531;
  reg [31:0] p23_add_64292;
  reg [31:0] p23_add_65634;
  reg [31:0] p23_add_64444;
  reg [31:0] p23_and_65715;
  reg [31:0] p23_add_65736;
  reg [31:0] p23_add_64445;
  reg [31:0] p23_add_64595;
  reg [31:0] p23_add_64480;
  reg [31:0] p23_add_64613;
  reg [31:0] p23_add_64631;
  reg [31:0] p23_add_64766;
  reg [31:0] p23_add_64904;
  reg [31:0] p23_add_65045;
  reg [31:0] p23_add_65186;
  reg [31:0] p23_add_65326;
  always_ff @ (posedge clk) begin
    p23_add_63929 <= p22_add_63929;
    p23_add_65503 <= p22_add_65503;
    p23_add_64256 <= p22_add_64256;
    p23_add_65607 <= p22_add_65607;
    p23_add_63999 <= p22_add_63999;
    p23_add_65707 <= p23_add_65707_comb;
    p23_add_65708 <= p23_add_65708_comb;
    p23_add_64275 <= p22_add_64275;
    p23_add_65714 <= p23_add_65714_comb;
    p23_add_65531 <= p22_add_65531;
    p23_add_64292 <= p22_add_64292;
    p23_add_65634 <= p22_add_65634;
    p23_add_64444 <= p22_add_64444;
    p23_and_65715 <= p23_and_65715_comb;
    p23_add_65736 <= p23_add_65736_comb;
    p23_add_64445 <= p22_add_64445;
    p23_add_64595 <= p22_add_64595;
    p23_add_64480 <= p22_add_64480;
    p23_add_64613 <= p22_add_64613;
    p23_add_64631 <= p22_add_64631;
    p23_add_64766 <= p22_add_64766;
    p23_add_64904 <= p22_add_64904;
    p23_add_65045 <= p22_add_65045;
    p23_add_65186 <= p22_add_65186;
    p23_add_65326 <= p22_add_65326;
  end

  // ===== Pipe stage 24:
  wire [31:0] p24_and_65817_comb;
  wire [31:0] p24_add_65808_comb;
  wire [30:0] p24_add_65813_comb;
  wire [31:0] p24_add_65809_comb;
  wire [31:0] p24_add_65836_comb;
  wire [31:0] p24_add_65810_comb;
  wire [31:0] p24_add_65816_comb;
  wire [31:0] p24_add_65838_comb;
  assign p24_and_65817_comb = p23_add_65736 & p23_add_65634;
  assign p24_add_65808_comb = (p23_add_65708 & p23_add_65607 ^ ~(p23_add_65708 | ~p23_add_65503)) + {p23_add_65708[5:0] ^ p23_add_65708[10:5] ^ p23_add_65708[24:19], p23_add_65708[31:27] ^ p23_add_65708[4:0] ^ p23_add_65708[18:14], p23_add_65708[26:13] ^ p23_add_65708[31:18] ^ p23_add_65708[13:0], p23_add_65708[12:6] ^ p23_add_65708[17:11] ^ p23_add_65708[31:25]};
  assign p24_add_65813_comb = p23_add_64292[31:1] + 31'h4c1f_28a9;
  assign p24_add_65809_comb = p24_add_65808_comb + p23_add_65714;
  assign p24_add_65836_comb = (p24_and_65817_comb ^ p23_add_65736 & p23_add_65531 ^ p23_and_65715) + p23_add_65707;
  assign p24_add_65810_comb = p24_add_65809_comb + p23_add_65531;
  assign p24_add_65816_comb = {p24_add_65813_comb, p23_add_64292[0]} + p23_add_65503;
  assign p24_add_65838_comb = p24_add_65836_comb + {p23_add_65736[1:0] ^ p23_add_65736[12:11] ^ p23_add_65736[21:20], p23_add_65736[31:21] ^ p23_add_65736[10:0] ^ p23_add_65736[19:9], p23_add_65736[20:12] ^ p23_add_65736[31:23] ^ p23_add_65736[8:0], p23_add_65736[11:2] ^ p23_add_65736[22:13] ^ p23_add_65736[31:22]};

  // Registers for pipe stage 24:
  reg [31:0] p24_add_63929;
  reg [31:0] p24_add_64256;
  reg [31:0] p24_add_65607;
  reg [31:0] p24_add_63999;
  reg [31:0] p24_add_65708;
  reg [31:0] p24_add_64275;
  reg [31:0] p24_add_65809;
  reg [31:0] p24_add_65810;
  reg [31:0] p24_add_64292;
  reg [31:0] p24_add_65816;
  reg [31:0] p24_add_65634;
  reg [31:0] p24_add_64444;
  reg [31:0] p24_add_65736;
  reg [31:0] p24_add_64445;
  reg [31:0] p24_and_65817;
  reg [31:0] p24_add_65838;
  reg [31:0] p24_add_64595;
  reg [31:0] p24_add_64480;
  reg [31:0] p24_add_64613;
  reg [31:0] p24_add_64631;
  reg [31:0] p24_add_64766;
  reg [31:0] p24_add_64904;
  reg [31:0] p24_add_65045;
  reg [31:0] p24_add_65186;
  reg [31:0] p24_add_65326;
  always_ff @ (posedge clk) begin
    p24_add_63929 <= p23_add_63929;
    p24_add_64256 <= p23_add_64256;
    p24_add_65607 <= p23_add_65607;
    p24_add_63999 <= p23_add_63999;
    p24_add_65708 <= p23_add_65708;
    p24_add_64275 <= p23_add_64275;
    p24_add_65809 <= p24_add_65809_comb;
    p24_add_65810 <= p24_add_65810_comb;
    p24_add_64292 <= p23_add_64292;
    p24_add_65816 <= p24_add_65816_comb;
    p24_add_65634 <= p23_add_65634;
    p24_add_64444 <= p23_add_64444;
    p24_add_65736 <= p23_add_65736;
    p24_add_64445 <= p23_add_64445;
    p24_and_65817 <= p24_and_65817_comb;
    p24_add_65838 <= p24_add_65838_comb;
    p24_add_64595 <= p23_add_64595;
    p24_add_64480 <= p23_add_64480;
    p24_add_64613 <= p23_add_64613;
    p24_add_64631 <= p23_add_64631;
    p24_add_64766 <= p23_add_64766;
    p24_add_64904 <= p23_add_64904;
    p24_add_65045 <= p23_add_65045;
    p24_add_65186 <= p23_add_65186;
    p24_add_65326 <= p23_add_65326;
  end

  // ===== Pipe stage 25:
  wire [31:0] p25_and_65916_comb;
  wire [31:0] p25_add_65910_comb;
  wire [31:0] p25_add_65911_comb;
  wire [31:0] p25_add_65914_comb;
  wire [31:0] p25_add_65935_comb;
  wire [31:0] p25_add_65912_comb;
  wire [31:0] p25_add_65915_comb;
  wire [31:0] p25_add_65937_comb;
  assign p25_and_65916_comb = p24_add_65838 & p24_add_65736;
  assign p25_add_65910_comb = (p24_add_65810 & p24_add_65708 ^ ~(p24_add_65810 | ~p24_add_65607)) + {p24_add_65810[5:0] ^ p24_add_65810[10:5] ^ p24_add_65810[24:19], p24_add_65810[31:27] ^ p24_add_65810[4:0] ^ p24_add_65810[18:14], p24_add_65810[26:13] ^ p24_add_65810[31:18] ^ p24_add_65810[13:0], p24_add_65810[12:6] ^ p24_add_65810[17:11] ^ p24_add_65810[31:25]};
  assign p25_add_65911_comb = p25_add_65910_comb + p24_add_65816;
  assign p25_add_65914_comb = p24_add_64444 + 32'ha831_c66d;
  assign p25_add_65935_comb = (p25_and_65916_comb ^ p24_add_65838 & p24_add_65634 ^ p24_and_65817) + p24_add_65809;
  assign p25_add_65912_comb = p25_add_65911_comb + p24_add_65634;
  assign p25_add_65915_comb = p24_add_65607 + p25_add_65914_comb;
  assign p25_add_65937_comb = p25_add_65935_comb + {p24_add_65838[1:0] ^ p24_add_65838[12:11] ^ p24_add_65838[21:20], p24_add_65838[31:21] ^ p24_add_65838[10:0] ^ p24_add_65838[19:9], p24_add_65838[20:12] ^ p24_add_65838[31:23] ^ p24_add_65838[8:0], p24_add_65838[11:2] ^ p24_add_65838[22:13] ^ p24_add_65838[31:22]};

  // Registers for pipe stage 25:
  reg [31:0] p25_add_63929;
  reg [31:0] p25_add_64256;
  reg [31:0] p25_add_63999;
  reg [31:0] p25_add_65708;
  reg [31:0] p25_add_64275;
  reg [31:0] p25_add_65810;
  reg [31:0] p25_add_64292;
  reg [31:0] p25_add_65911;
  reg [31:0] p25_add_65912;
  reg [31:0] p25_add_64444;
  reg [31:0] p25_add_65915;
  reg [31:0] p25_add_65736;
  reg [31:0] p25_add_64445;
  reg [31:0] p25_add_65838;
  reg [31:0] p25_add_64595;
  reg [31:0] p25_and_65916;
  reg [31:0] p25_add_65937;
  reg [31:0] p25_add_64480;
  reg [31:0] p25_add_64613;
  reg [31:0] p25_add_64631;
  reg [31:0] p25_add_64766;
  reg [31:0] p25_add_64904;
  reg [31:0] p25_add_65045;
  reg [31:0] p25_add_65186;
  reg [31:0] p25_add_65326;
  always_ff @ (posedge clk) begin
    p25_add_63929 <= p24_add_63929;
    p25_add_64256 <= p24_add_64256;
    p25_add_63999 <= p24_add_63999;
    p25_add_65708 <= p24_add_65708;
    p25_add_64275 <= p24_add_64275;
    p25_add_65810 <= p24_add_65810;
    p25_add_64292 <= p24_add_64292;
    p25_add_65911 <= p25_add_65911_comb;
    p25_add_65912 <= p25_add_65912_comb;
    p25_add_64444 <= p24_add_64444;
    p25_add_65915 <= p25_add_65915_comb;
    p25_add_65736 <= p24_add_65736;
    p25_add_64445 <= p24_add_64445;
    p25_add_65838 <= p24_add_65838;
    p25_add_64595 <= p24_add_64595;
    p25_and_65916 <= p25_and_65916_comb;
    p25_add_65937 <= p25_add_65937_comb;
    p25_add_64480 <= p24_add_64480;
    p25_add_64613 <= p24_add_64613;
    p25_add_64631 <= p24_add_64631;
    p25_add_64766 <= p24_add_64766;
    p25_add_64904 <= p24_add_64904;
    p25_add_65045 <= p24_add_65045;
    p25_add_65186 <= p24_add_65186;
    p25_add_65326 <= p24_add_65326;
  end

  // ===== Pipe stage 26:
  wire [31:0] p26_and_66018_comb;
  wire [31:0] p26_add_66009_comb;
  wire [28:0] p26_add_66014_comb;
  wire [31:0] p26_add_66010_comb;
  wire [31:0] p26_add_66037_comb;
  wire [31:0] p26_add_66011_comb;
  wire [31:0] p26_add_66017_comb;
  wire [31:0] p26_add_66039_comb;
  assign p26_and_66018_comb = p25_add_65937 & p25_add_65838;
  assign p26_add_66009_comb = {p25_add_65912[5:0] ^ p25_add_65912[10:5] ^ p25_add_65912[24:19], p25_add_65912[31:27] ^ p25_add_65912[4:0] ^ p25_add_65912[18:14], p25_add_65912[26:13] ^ p25_add_65912[31:18] ^ p25_add_65912[13:0], p25_add_65912[12:6] ^ p25_add_65912[17:11] ^ p25_add_65912[31:25]} + (p25_add_65912 & p25_add_65810 ^ ~(p25_add_65912 | ~p25_add_65708));
  assign p26_add_66014_comb = p25_add_64445[31:3] + 29'h1600_64f9;
  assign p26_add_66010_comb = p26_add_66009_comb + p25_add_65915;
  assign p26_add_66037_comb = (p26_and_66018_comb ^ p25_add_65937 & p25_add_65736 ^ p25_and_65916) + p25_add_65911;
  assign p26_add_66011_comb = p26_add_66010_comb + p25_add_65736;
  assign p26_add_66017_comb = {p26_add_66014_comb, p25_add_64445[2:0]} + p25_add_65708;
  assign p26_add_66039_comb = p26_add_66037_comb + {p25_add_65937[1:0] ^ p25_add_65937[12:11] ^ p25_add_65937[21:20], p25_add_65937[31:21] ^ p25_add_65937[10:0] ^ p25_add_65937[19:9], p25_add_65937[20:12] ^ p25_add_65937[31:23] ^ p25_add_65937[8:0], p25_add_65937[11:2] ^ p25_add_65937[22:13] ^ p25_add_65937[31:22]};

  // Registers for pipe stage 26:
  reg [31:0] p26_add_63929;
  reg [31:0] p26_add_64256;
  reg [31:0] p26_add_63999;
  reg [31:0] p26_add_64275;
  reg [31:0] p26_add_65810;
  reg [31:0] p26_add_64292;
  reg [31:0] p26_add_65912;
  reg [31:0] p26_add_64444;
  reg [31:0] p26_add_66010;
  reg [31:0] p26_add_66011;
  reg [31:0] p26_add_64445;
  reg [31:0] p26_add_66017;
  reg [31:0] p26_add_65838;
  reg [31:0] p26_add_64595;
  reg [31:0] p26_add_65937;
  reg [31:0] p26_add_64480;
  reg [31:0] p26_and_66018;
  reg [31:0] p26_add_66039;
  reg [31:0] p26_add_64613;
  reg [31:0] p26_add_64631;
  reg [31:0] p26_add_64766;
  reg [31:0] p26_add_64904;
  reg [31:0] p26_add_65045;
  reg [31:0] p26_add_65186;
  reg [31:0] p26_add_65326;
  always_ff @ (posedge clk) begin
    p26_add_63929 <= p25_add_63929;
    p26_add_64256 <= p25_add_64256;
    p26_add_63999 <= p25_add_63999;
    p26_add_64275 <= p25_add_64275;
    p26_add_65810 <= p25_add_65810;
    p26_add_64292 <= p25_add_64292;
    p26_add_65912 <= p25_add_65912;
    p26_add_64444 <= p25_add_64444;
    p26_add_66010 <= p26_add_66010_comb;
    p26_add_66011 <= p26_add_66011_comb;
    p26_add_64445 <= p25_add_64445;
    p26_add_66017 <= p26_add_66017_comb;
    p26_add_65838 <= p25_add_65838;
    p26_add_64595 <= p25_add_64595;
    p26_add_65937 <= p25_add_65937;
    p26_add_64480 <= p25_add_64480;
    p26_and_66018 <= p26_and_66018_comb;
    p26_add_66039 <= p26_add_66039_comb;
    p26_add_64613 <= p25_add_64613;
    p26_add_64631 <= p25_add_64631;
    p26_add_64766 <= p25_add_64766;
    p26_add_64904 <= p25_add_64904;
    p26_add_65045 <= p25_add_65045;
    p26_add_65186 <= p25_add_65186;
    p26_add_65326 <= p25_add_65326;
  end

  // ===== Pipe stage 27:
  wire [31:0] p27_and_66117_comb;
  wire [31:0] p27_add_66111_comb;
  wire [31:0] p27_add_66112_comb;
  wire [31:0] p27_add_66115_comb;
  wire [31:0] p27_add_66136_comb;
  wire [31:0] p27_add_66113_comb;
  wire [31:0] p27_add_66116_comb;
  wire [31:0] p27_add_66138_comb;
  assign p27_and_66117_comb = p26_add_66039 & p26_add_65937;
  assign p27_add_66111_comb = (p26_add_66011 & p26_add_65912 ^ ~(p26_add_66011 | ~p26_add_65810)) + {p26_add_66011[5:0] ^ p26_add_66011[10:5] ^ p26_add_66011[24:19], p26_add_66011[31:27] ^ p26_add_66011[4:0] ^ p26_add_66011[18:14], p26_add_66011[26:13] ^ p26_add_66011[31:18] ^ p26_add_66011[13:0], p26_add_66011[12:6] ^ p26_add_66011[17:11] ^ p26_add_66011[31:25]};
  assign p27_add_66112_comb = p27_add_66111_comb + p26_add_66017;
  assign p27_add_66115_comb = p26_add_64595 + 32'hbf59_7fc7;
  assign p27_add_66136_comb = (p27_and_66117_comb ^ p26_add_66039 & p26_add_65838 ^ p26_and_66018) + p26_add_66010;
  assign p27_add_66113_comb = p27_add_66112_comb + p26_add_65838;
  assign p27_add_66116_comb = p26_add_65810 + p27_add_66115_comb;
  assign p27_add_66138_comb = p27_add_66136_comb + {p26_add_66039[1:0] ^ p26_add_66039[12:11] ^ p26_add_66039[21:20], p26_add_66039[31:21] ^ p26_add_66039[10:0] ^ p26_add_66039[19:9], p26_add_66039[20:12] ^ p26_add_66039[31:23] ^ p26_add_66039[8:0], p26_add_66039[11:2] ^ p26_add_66039[22:13] ^ p26_add_66039[31:22]};

  // Registers for pipe stage 27:
  reg [31:0] p27_add_63929;
  reg [31:0] p27_add_64256;
  reg [31:0] p27_add_63999;
  reg [31:0] p27_add_64275;
  reg [31:0] p27_add_64292;
  reg [31:0] p27_add_65912;
  reg [31:0] p27_add_64444;
  reg [31:0] p27_add_66011;
  reg [31:0] p27_add_64445;
  reg [31:0] p27_add_66112;
  reg [31:0] p27_add_66113;
  reg [31:0] p27_add_64595;
  reg [31:0] p27_add_66116;
  reg [31:0] p27_add_65937;
  reg [31:0] p27_add_64480;
  reg [31:0] p27_add_66039;
  reg [31:0] p27_add_64613;
  reg [31:0] p27_and_66117;
  reg [31:0] p27_add_66138;
  reg [31:0] p27_add_64631;
  reg [31:0] p27_add_64766;
  reg [31:0] p27_add_64904;
  reg [31:0] p27_add_65045;
  reg [31:0] p27_add_65186;
  reg [31:0] p27_add_65326;
  always_ff @ (posedge clk) begin
    p27_add_63929 <= p26_add_63929;
    p27_add_64256 <= p26_add_64256;
    p27_add_63999 <= p26_add_63999;
    p27_add_64275 <= p26_add_64275;
    p27_add_64292 <= p26_add_64292;
    p27_add_65912 <= p26_add_65912;
    p27_add_64444 <= p26_add_64444;
    p27_add_66011 <= p26_add_66011;
    p27_add_64445 <= p26_add_64445;
    p27_add_66112 <= p27_add_66112_comb;
    p27_add_66113 <= p27_add_66113_comb;
    p27_add_64595 <= p26_add_64595;
    p27_add_66116 <= p27_add_66116_comb;
    p27_add_65937 <= p26_add_65937;
    p27_add_64480 <= p26_add_64480;
    p27_add_66039 <= p26_add_66039;
    p27_add_64613 <= p26_add_64613;
    p27_and_66117 <= p27_and_66117_comb;
    p27_add_66138 <= p27_add_66138_comb;
    p27_add_64631 <= p26_add_64631;
    p27_add_64766 <= p26_add_64766;
    p27_add_64904 <= p26_add_64904;
    p27_add_65045 <= p26_add_65045;
    p27_add_65186 <= p26_add_65186;
    p27_add_65326 <= p26_add_65326;
  end

  // ===== Pipe stage 28:
  wire [31:0] p28_and_66216_comb;
  wire [31:0] p28_add_66210_comb;
  wire [31:0] p28_add_66211_comb;
  wire [31:0] p28_add_66214_comb;
  wire [31:0] p28_add_66235_comb;
  wire [31:0] p28_add_66212_comb;
  wire [31:0] p28_add_66215_comb;
  wire [31:0] p28_add_66237_comb;
  assign p28_and_66216_comb = p27_add_66138 & p27_add_66039;
  assign p28_add_66210_comb = {p27_add_66113[5:0] ^ p27_add_66113[10:5] ^ p27_add_66113[24:19], p27_add_66113[31:27] ^ p27_add_66113[4:0] ^ p27_add_66113[18:14], p27_add_66113[26:13] ^ p27_add_66113[31:18] ^ p27_add_66113[13:0], p27_add_66113[12:6] ^ p27_add_66113[17:11] ^ p27_add_66113[31:25]} + (p27_add_66113 & p27_add_66011 ^ ~(p27_add_66113 | ~p27_add_65912));
  assign p28_add_66211_comb = p28_add_66210_comb + p27_add_66116;
  assign p28_add_66214_comb = p27_add_64480 + 32'hc6e0_0bf3;
  assign p28_add_66235_comb = (p28_and_66216_comb ^ p27_add_66138 & p27_add_65937 ^ p27_and_66117) + p27_add_66112;
  assign p28_add_66212_comb = p28_add_66211_comb + p27_add_65937;
  assign p28_add_66215_comb = p27_add_65912 + p28_add_66214_comb;
  assign p28_add_66237_comb = p28_add_66235_comb + {p27_add_66138[1:0] ^ p27_add_66138[12:11] ^ p27_add_66138[21:20], p27_add_66138[31:21] ^ p27_add_66138[10:0] ^ p27_add_66138[19:9], p27_add_66138[20:12] ^ p27_add_66138[31:23] ^ p27_add_66138[8:0], p27_add_66138[11:2] ^ p27_add_66138[22:13] ^ p27_add_66138[31:22]};

  // Registers for pipe stage 28:
  reg [31:0] p28_add_63929;
  reg [31:0] p28_add_64256;
  reg [31:0] p28_add_63999;
  reg [31:0] p28_add_64275;
  reg [31:0] p28_add_64292;
  reg [31:0] p28_add_64444;
  reg [31:0] p28_add_66011;
  reg [31:0] p28_add_64445;
  reg [31:0] p28_add_66113;
  reg [31:0] p28_add_64595;
  reg [31:0] p28_add_66211;
  reg [31:0] p28_add_66212;
  reg [31:0] p28_add_64480;
  reg [31:0] p28_add_66215;
  reg [31:0] p28_add_66039;
  reg [31:0] p28_add_64613;
  reg [31:0] p28_add_66138;
  reg [31:0] p28_add_64631;
  reg [31:0] p28_and_66216;
  reg [31:0] p28_add_66237;
  reg [31:0] p28_add_64766;
  reg [31:0] p28_add_64904;
  reg [31:0] p28_add_65045;
  reg [31:0] p28_add_65186;
  reg [31:0] p28_add_65326;
  always_ff @ (posedge clk) begin
    p28_add_63929 <= p27_add_63929;
    p28_add_64256 <= p27_add_64256;
    p28_add_63999 <= p27_add_63999;
    p28_add_64275 <= p27_add_64275;
    p28_add_64292 <= p27_add_64292;
    p28_add_64444 <= p27_add_64444;
    p28_add_66011 <= p27_add_66011;
    p28_add_64445 <= p27_add_64445;
    p28_add_66113 <= p27_add_66113;
    p28_add_64595 <= p27_add_64595;
    p28_add_66211 <= p28_add_66211_comb;
    p28_add_66212 <= p28_add_66212_comb;
    p28_add_64480 <= p27_add_64480;
    p28_add_66215 <= p28_add_66215_comb;
    p28_add_66039 <= p27_add_66039;
    p28_add_64613 <= p27_add_64613;
    p28_add_66138 <= p27_add_66138;
    p28_add_64631 <= p27_add_64631;
    p28_and_66216 <= p28_and_66216_comb;
    p28_add_66237 <= p28_add_66237_comb;
    p28_add_64766 <= p27_add_64766;
    p28_add_64904 <= p27_add_64904;
    p28_add_65045 <= p27_add_65045;
    p28_add_65186 <= p27_add_65186;
    p28_add_65326 <= p27_add_65326;
  end

  // ===== Pipe stage 29:
  wire [31:0] p29_and_66315_comb;
  wire [31:0] p29_add_66309_comb;
  wire [31:0] p29_add_66310_comb;
  wire [31:0] p29_add_66313_comb;
  wire [31:0] p29_add_66334_comb;
  wire [31:0] p29_add_66311_comb;
  wire [31:0] p29_add_66314_comb;
  wire [31:0] p29_add_66336_comb;
  assign p29_and_66315_comb = p28_add_66237 & p28_add_66138;
  assign p29_add_66309_comb = {p28_add_66212[5:0] ^ p28_add_66212[10:5] ^ p28_add_66212[24:19], p28_add_66212[31:27] ^ p28_add_66212[4:0] ^ p28_add_66212[18:14], p28_add_66212[26:13] ^ p28_add_66212[31:18] ^ p28_add_66212[13:0], p28_add_66212[12:6] ^ p28_add_66212[17:11] ^ p28_add_66212[31:25]} + (p28_add_66212 & p28_add_66113 ^ ~(p28_add_66212 | ~p28_add_66011));
  assign p29_add_66310_comb = p29_add_66309_comb + p28_add_66215;
  assign p29_add_66313_comb = p28_add_64613 + 32'hd5a7_9147;
  assign p29_add_66334_comb = (p29_and_66315_comb ^ p28_add_66237 & p28_add_66039 ^ p28_and_66216) + p28_add_66211;
  assign p29_add_66311_comb = p29_add_66310_comb + p28_add_66039;
  assign p29_add_66314_comb = p28_add_66011 + p29_add_66313_comb;
  assign p29_add_66336_comb = p29_add_66334_comb + {p28_add_66237[1:0] ^ p28_add_66237[12:11] ^ p28_add_66237[21:20], p28_add_66237[31:21] ^ p28_add_66237[10:0] ^ p28_add_66237[19:9], p28_add_66237[20:12] ^ p28_add_66237[31:23] ^ p28_add_66237[8:0], p28_add_66237[11:2] ^ p28_add_66237[22:13] ^ p28_add_66237[31:22]};

  // Registers for pipe stage 29:
  reg [31:0] p29_add_63929;
  reg [31:0] p29_add_64256;
  reg [31:0] p29_add_63999;
  reg [31:0] p29_add_64275;
  reg [31:0] p29_add_64292;
  reg [31:0] p29_add_64444;
  reg [31:0] p29_add_64445;
  reg [31:0] p29_add_66113;
  reg [31:0] p29_add_64595;
  reg [31:0] p29_add_66212;
  reg [31:0] p29_add_64480;
  reg [31:0] p29_add_66310;
  reg [31:0] p29_add_66311;
  reg [31:0] p29_add_64613;
  reg [31:0] p29_add_66314;
  reg [31:0] p29_add_66138;
  reg [31:0] p29_add_64631;
  reg [31:0] p29_add_66237;
  reg [31:0] p29_add_64766;
  reg [31:0] p29_and_66315;
  reg [31:0] p29_add_66336;
  reg [31:0] p29_add_64904;
  reg [31:0] p29_add_65045;
  reg [31:0] p29_add_65186;
  reg [31:0] p29_add_65326;
  always_ff @ (posedge clk) begin
    p29_add_63929 <= p28_add_63929;
    p29_add_64256 <= p28_add_64256;
    p29_add_63999 <= p28_add_63999;
    p29_add_64275 <= p28_add_64275;
    p29_add_64292 <= p28_add_64292;
    p29_add_64444 <= p28_add_64444;
    p29_add_64445 <= p28_add_64445;
    p29_add_66113 <= p28_add_66113;
    p29_add_64595 <= p28_add_64595;
    p29_add_66212 <= p28_add_66212;
    p29_add_64480 <= p28_add_64480;
    p29_add_66310 <= p29_add_66310_comb;
    p29_add_66311 <= p29_add_66311_comb;
    p29_add_64613 <= p28_add_64613;
    p29_add_66314 <= p29_add_66314_comb;
    p29_add_66138 <= p28_add_66138;
    p29_add_64631 <= p28_add_64631;
    p29_add_66237 <= p28_add_66237;
    p29_add_64766 <= p28_add_64766;
    p29_and_66315 <= p29_and_66315_comb;
    p29_add_66336 <= p29_add_66336_comb;
    p29_add_64904 <= p28_add_64904;
    p29_add_65045 <= p28_add_65045;
    p29_add_65186 <= p28_add_65186;
    p29_add_65326 <= p28_add_65326;
  end

  // ===== Pipe stage 30:
  wire [31:0] p30_and_66414_comb;
  wire [31:0] p30_add_66408_comb;
  wire [31:0] p30_add_66409_comb;
  wire [31:0] p30_add_66412_comb;
  wire [31:0] p30_add_66433_comb;
  wire [31:0] p30_add_66410_comb;
  wire [31:0] p30_add_66413_comb;
  wire [31:0] p30_add_66435_comb;
  assign p30_and_66414_comb = p29_add_66336 & p29_add_66237;
  assign p30_add_66408_comb = {p29_add_66311[5:0] ^ p29_add_66311[10:5] ^ p29_add_66311[24:19], p29_add_66311[31:27] ^ p29_add_66311[4:0] ^ p29_add_66311[18:14], p29_add_66311[26:13] ^ p29_add_66311[31:18] ^ p29_add_66311[13:0], p29_add_66311[12:6] ^ p29_add_66311[17:11] ^ p29_add_66311[31:25]} + (p29_add_66311 & p29_add_66212 ^ ~(p29_add_66311 | ~p29_add_66113));
  assign p30_add_66409_comb = p30_add_66408_comb + p29_add_66314;
  assign p30_add_66412_comb = p29_add_64631 + 32'h06ca_6351;
  assign p30_add_66433_comb = (p30_and_66414_comb ^ p29_add_66336 & p29_add_66138 ^ p29_and_66315) + p29_add_66310;
  assign p30_add_66410_comb = p30_add_66409_comb + p29_add_66138;
  assign p30_add_66413_comb = p29_add_66113 + p30_add_66412_comb;
  assign p30_add_66435_comb = p30_add_66433_comb + {p29_add_66336[1:0] ^ p29_add_66336[12:11] ^ p29_add_66336[21:20], p29_add_66336[31:21] ^ p29_add_66336[10:0] ^ p29_add_66336[19:9], p29_add_66336[20:12] ^ p29_add_66336[31:23] ^ p29_add_66336[8:0], p29_add_66336[11:2] ^ p29_add_66336[22:13] ^ p29_add_66336[31:22]};

  // Registers for pipe stage 30:
  reg [31:0] p30_add_63929;
  reg [31:0] p30_add_64256;
  reg [31:0] p30_add_63999;
  reg [31:0] p30_add_64275;
  reg [31:0] p30_add_64292;
  reg [31:0] p30_add_64444;
  reg [31:0] p30_add_64445;
  reg [31:0] p30_add_64595;
  reg [31:0] p30_add_66212;
  reg [31:0] p30_add_64480;
  reg [31:0] p30_add_66311;
  reg [31:0] p30_add_64613;
  reg [31:0] p30_add_66409;
  reg [31:0] p30_add_66410;
  reg [31:0] p30_add_64631;
  reg [31:0] p30_add_66413;
  reg [31:0] p30_add_66237;
  reg [31:0] p30_add_64766;
  reg [31:0] p30_add_66336;
  reg [31:0] p30_add_64904;
  reg [31:0] p30_and_66414;
  reg [31:0] p30_add_66435;
  reg [31:0] p30_add_65045;
  reg [31:0] p30_add_65186;
  reg [31:0] p30_add_65326;
  always_ff @ (posedge clk) begin
    p30_add_63929 <= p29_add_63929;
    p30_add_64256 <= p29_add_64256;
    p30_add_63999 <= p29_add_63999;
    p30_add_64275 <= p29_add_64275;
    p30_add_64292 <= p29_add_64292;
    p30_add_64444 <= p29_add_64444;
    p30_add_64445 <= p29_add_64445;
    p30_add_64595 <= p29_add_64595;
    p30_add_66212 <= p29_add_66212;
    p30_add_64480 <= p29_add_64480;
    p30_add_66311 <= p29_add_66311;
    p30_add_64613 <= p29_add_64613;
    p30_add_66409 <= p30_add_66409_comb;
    p30_add_66410 <= p30_add_66410_comb;
    p30_add_64631 <= p29_add_64631;
    p30_add_66413 <= p30_add_66413_comb;
    p30_add_66237 <= p29_add_66237;
    p30_add_64766 <= p29_add_64766;
    p30_add_66336 <= p29_add_66336;
    p30_add_64904 <= p29_add_64904;
    p30_and_66414 <= p30_and_66414_comb;
    p30_add_66435 <= p30_add_66435_comb;
    p30_add_65045 <= p29_add_65045;
    p30_add_65186 <= p29_add_65186;
    p30_add_65326 <= p29_add_65326;
  end

  // ===== Pipe stage 31:
  wire [31:0] p31_and_66513_comb;
  wire [31:0] p31_add_66507_comb;
  wire [31:0] p31_add_66508_comb;
  wire [31:0] p31_add_66511_comb;
  wire [31:0] p31_add_66532_comb;
  wire [31:0] p31_add_66509_comb;
  wire [31:0] p31_add_66512_comb;
  wire [31:0] p31_add_66534_comb;
  assign p31_and_66513_comb = p30_add_66435 & p30_add_66336;
  assign p31_add_66507_comb = {p30_add_66410[5:0] ^ p30_add_66410[10:5] ^ p30_add_66410[24:19], p30_add_66410[31:27] ^ p30_add_66410[4:0] ^ p30_add_66410[18:14], p30_add_66410[26:13] ^ p30_add_66410[31:18] ^ p30_add_66410[13:0], p30_add_66410[12:6] ^ p30_add_66410[17:11] ^ p30_add_66410[31:25]} + (p30_add_66410 & p30_add_66311 ^ ~(p30_add_66410 | ~p30_add_66212));
  assign p31_add_66508_comb = p31_add_66507_comb + p30_add_66413;
  assign p31_add_66511_comb = p30_add_64766 + 32'h1429_2967;
  assign p31_add_66532_comb = (p31_and_66513_comb ^ p30_add_66435 & p30_add_66237 ^ p30_and_66414) + p30_add_66409;
  assign p31_add_66509_comb = p31_add_66508_comb + p30_add_66237;
  assign p31_add_66512_comb = p30_add_66212 + p31_add_66511_comb;
  assign p31_add_66534_comb = p31_add_66532_comb + {p30_add_66435[1:0] ^ p30_add_66435[12:11] ^ p30_add_66435[21:20], p30_add_66435[31:21] ^ p30_add_66435[10:0] ^ p30_add_66435[19:9], p30_add_66435[20:12] ^ p30_add_66435[31:23] ^ p30_add_66435[8:0], p30_add_66435[11:2] ^ p30_add_66435[22:13] ^ p30_add_66435[31:22]};

  // Registers for pipe stage 31:
  reg [31:0] p31_add_63929;
  reg [31:0] p31_add_64256;
  reg [31:0] p31_add_63999;
  reg [31:0] p31_add_64275;
  reg [31:0] p31_add_64292;
  reg [31:0] p31_add_64444;
  reg [31:0] p31_add_64445;
  reg [31:0] p31_add_64595;
  reg [31:0] p31_add_64480;
  reg [31:0] p31_add_66311;
  reg [31:0] p31_add_64613;
  reg [31:0] p31_add_66410;
  reg [31:0] p31_add_64631;
  reg [31:0] p31_add_66508;
  reg [31:0] p31_add_66509;
  reg [31:0] p31_add_64766;
  reg [31:0] p31_add_66512;
  reg [31:0] p31_add_66336;
  reg [31:0] p31_add_64904;
  reg [31:0] p31_add_66435;
  reg [31:0] p31_add_65045;
  reg [31:0] p31_and_66513;
  reg [31:0] p31_add_66534;
  reg [31:0] p31_add_65186;
  reg [31:0] p31_add_65326;
  always_ff @ (posedge clk) begin
    p31_add_63929 <= p30_add_63929;
    p31_add_64256 <= p30_add_64256;
    p31_add_63999 <= p30_add_63999;
    p31_add_64275 <= p30_add_64275;
    p31_add_64292 <= p30_add_64292;
    p31_add_64444 <= p30_add_64444;
    p31_add_64445 <= p30_add_64445;
    p31_add_64595 <= p30_add_64595;
    p31_add_64480 <= p30_add_64480;
    p31_add_66311 <= p30_add_66311;
    p31_add_64613 <= p30_add_64613;
    p31_add_66410 <= p30_add_66410;
    p31_add_64631 <= p30_add_64631;
    p31_add_66508 <= p31_add_66508_comb;
    p31_add_66509 <= p31_add_66509_comb;
    p31_add_64766 <= p30_add_64766;
    p31_add_66512 <= p31_add_66512_comb;
    p31_add_66336 <= p30_add_66336;
    p31_add_64904 <= p30_add_64904;
    p31_add_66435 <= p30_add_66435;
    p31_add_65045 <= p30_add_65045;
    p31_and_66513 <= p31_and_66513_comb;
    p31_add_66534 <= p31_add_66534_comb;
    p31_add_65186 <= p30_add_65186;
    p31_add_65326 <= p30_add_65326;
  end

  // ===== Pipe stage 32:
  wire [31:0] p32_and_66612_comb;
  wire [31:0] p32_add_66606_comb;
  wire [31:0] p32_add_66607_comb;
  wire [31:0] p32_add_66610_comb;
  wire [31:0] p32_add_66631_comb;
  wire [31:0] p32_add_66608_comb;
  wire [31:0] p32_add_66611_comb;
  wire [31:0] p32_add_66633_comb;
  assign p32_and_66612_comb = p31_add_66534 & p31_add_66435;
  assign p32_add_66606_comb = {p31_add_66509[5:0] ^ p31_add_66509[10:5] ^ p31_add_66509[24:19], p31_add_66509[31:27] ^ p31_add_66509[4:0] ^ p31_add_66509[18:14], p31_add_66509[26:13] ^ p31_add_66509[31:18] ^ p31_add_66509[13:0], p31_add_66509[12:6] ^ p31_add_66509[17:11] ^ p31_add_66509[31:25]} + (p31_add_66509 & p31_add_66410 ^ ~(p31_add_66509 | ~p31_add_66311));
  assign p32_add_66607_comb = p32_add_66606_comb + p31_add_66512;
  assign p32_add_66610_comb = p31_add_64904 + 32'h27b7_0a85;
  assign p32_add_66631_comb = (p32_and_66612_comb ^ p31_add_66534 & p31_add_66336 ^ p31_and_66513) + p31_add_66508;
  assign p32_add_66608_comb = p32_add_66607_comb + p31_add_66336;
  assign p32_add_66611_comb = p31_add_66311 + p32_add_66610_comb;
  assign p32_add_66633_comb = p32_add_66631_comb + {p31_add_66534[1:0] ^ p31_add_66534[12:11] ^ p31_add_66534[21:20], p31_add_66534[31:21] ^ p31_add_66534[10:0] ^ p31_add_66534[19:9], p31_add_66534[20:12] ^ p31_add_66534[31:23] ^ p31_add_66534[8:0], p31_add_66534[11:2] ^ p31_add_66534[22:13] ^ p31_add_66534[31:22]};

  // Registers for pipe stage 32:
  reg [31:0] p32_add_63929;
  reg [31:0] p32_add_64256;
  reg [31:0] p32_add_63999;
  reg [31:0] p32_add_64275;
  reg [31:0] p32_add_64292;
  reg [31:0] p32_add_64444;
  reg [31:0] p32_add_64445;
  reg [31:0] p32_add_64595;
  reg [31:0] p32_add_64480;
  reg [31:0] p32_add_64613;
  reg [31:0] p32_add_66410;
  reg [31:0] p32_add_64631;
  reg [31:0] p32_add_66509;
  reg [31:0] p32_add_64766;
  reg [31:0] p32_add_66607;
  reg [31:0] p32_add_66608;
  reg [31:0] p32_add_64904;
  reg [31:0] p32_add_66611;
  reg [31:0] p32_add_66435;
  reg [31:0] p32_add_65045;
  reg [31:0] p32_add_66534;
  reg [31:0] p32_add_65186;
  reg [31:0] p32_and_66612;
  reg [31:0] p32_add_66633;
  reg [31:0] p32_add_65326;
  always_ff @ (posedge clk) begin
    p32_add_63929 <= p31_add_63929;
    p32_add_64256 <= p31_add_64256;
    p32_add_63999 <= p31_add_63999;
    p32_add_64275 <= p31_add_64275;
    p32_add_64292 <= p31_add_64292;
    p32_add_64444 <= p31_add_64444;
    p32_add_64445 <= p31_add_64445;
    p32_add_64595 <= p31_add_64595;
    p32_add_64480 <= p31_add_64480;
    p32_add_64613 <= p31_add_64613;
    p32_add_66410 <= p31_add_66410;
    p32_add_64631 <= p31_add_64631;
    p32_add_66509 <= p31_add_66509;
    p32_add_64766 <= p31_add_64766;
    p32_add_66607 <= p32_add_66607_comb;
    p32_add_66608 <= p32_add_66608_comb;
    p32_add_64904 <= p31_add_64904;
    p32_add_66611 <= p32_add_66611_comb;
    p32_add_66435 <= p31_add_66435;
    p32_add_65045 <= p31_add_65045;
    p32_add_66534 <= p31_add_66534;
    p32_add_65186 <= p31_add_65186;
    p32_and_66612 <= p32_and_66612_comb;
    p32_add_66633 <= p32_add_66633_comb;
    p32_add_65326 <= p31_add_65326;
  end

  // ===== Pipe stage 33:
  wire [31:0] p33_and_66714_comb;
  wire [31:0] p33_add_66705_comb;
  wire [28:0] p33_add_66710_comb;
  wire [31:0] p33_add_66706_comb;
  wire [31:0] p33_add_66733_comb;
  wire [31:0] p33_add_66707_comb;
  wire [31:0] p33_add_66713_comb;
  wire [31:0] p33_add_66735_comb;
  assign p33_and_66714_comb = p32_add_66633 & p32_add_66534;
  assign p33_add_66705_comb = {p32_add_66608[5:0] ^ p32_add_66608[10:5] ^ p32_add_66608[24:19], p32_add_66608[31:27] ^ p32_add_66608[4:0] ^ p32_add_66608[18:14], p32_add_66608[26:13] ^ p32_add_66608[31:18] ^ p32_add_66608[13:0], p32_add_66608[12:6] ^ p32_add_66608[17:11] ^ p32_add_66608[31:25]} + (p32_add_66608 & p32_add_66509 ^ ~(p32_add_66608 | ~p32_add_66410));
  assign p33_add_66710_comb = p32_add_65045[31:3] + 29'h05c3_6427;
  assign p33_add_66706_comb = p33_add_66705_comb + p32_add_66611;
  assign p33_add_66733_comb = (p33_and_66714_comb ^ p32_add_66633 & p32_add_66435 ^ p32_and_66612) + p32_add_66607;
  assign p33_add_66707_comb = p33_add_66706_comb + p32_add_66435;
  assign p33_add_66713_comb = {p33_add_66710_comb, p32_add_65045[2:0]} + p32_add_66410;
  assign p33_add_66735_comb = p33_add_66733_comb + {p32_add_66633[1:0] ^ p32_add_66633[12:11] ^ p32_add_66633[21:20], p32_add_66633[31:21] ^ p32_add_66633[10:0] ^ p32_add_66633[19:9], p32_add_66633[20:12] ^ p32_add_66633[31:23] ^ p32_add_66633[8:0], p32_add_66633[11:2] ^ p32_add_66633[22:13] ^ p32_add_66633[31:22]};

  // Registers for pipe stage 33:
  reg [31:0] p33_add_63929;
  reg [31:0] p33_add_64256;
  reg [31:0] p33_add_63999;
  reg [31:0] p33_add_64275;
  reg [31:0] p33_add_64292;
  reg [31:0] p33_add_64444;
  reg [31:0] p33_add_64445;
  reg [31:0] p33_add_64595;
  reg [31:0] p33_add_64480;
  reg [31:0] p33_add_64613;
  reg [31:0] p33_add_64631;
  reg [31:0] p33_add_66509;
  reg [31:0] p33_add_64766;
  reg [31:0] p33_add_66608;
  reg [31:0] p33_add_64904;
  reg [31:0] p33_add_66706;
  reg [31:0] p33_add_66707;
  reg [31:0] p33_add_65045;
  reg [31:0] p33_add_66713;
  reg [31:0] p33_add_66534;
  reg [31:0] p33_add_65186;
  reg [31:0] p33_add_66633;
  reg [31:0] p33_add_65326;
  reg [31:0] p33_and_66714;
  reg [31:0] p33_add_66735;
  always_ff @ (posedge clk) begin
    p33_add_63929 <= p32_add_63929;
    p33_add_64256 <= p32_add_64256;
    p33_add_63999 <= p32_add_63999;
    p33_add_64275 <= p32_add_64275;
    p33_add_64292 <= p32_add_64292;
    p33_add_64444 <= p32_add_64444;
    p33_add_64445 <= p32_add_64445;
    p33_add_64595 <= p32_add_64595;
    p33_add_64480 <= p32_add_64480;
    p33_add_64613 <= p32_add_64613;
    p33_add_64631 <= p32_add_64631;
    p33_add_66509 <= p32_add_66509;
    p33_add_64766 <= p32_add_64766;
    p33_add_66608 <= p32_add_66608;
    p33_add_64904 <= p32_add_64904;
    p33_add_66706 <= p33_add_66706_comb;
    p33_add_66707 <= p33_add_66707_comb;
    p33_add_65045 <= p32_add_65045;
    p33_add_66713 <= p33_add_66713_comb;
    p33_add_66534 <= p32_add_66534;
    p33_add_65186 <= p32_add_65186;
    p33_add_66633 <= p32_add_66633;
    p33_add_65326 <= p32_add_65326;
    p33_and_66714 <= p33_and_66714_comb;
    p33_add_66735 <= p33_add_66735_comb;
  end

  // ===== Pipe stage 34:
  wire [31:0] p34_and_66850_comb;
  wire [31:0] p34_add_66807_comb;
  wire [29:0] p34_add_66812_comb;
  wire [31:0] p34_add_66808_comb;
  wire [31:0] p34_add_66847_comb;
  wire [31:0] p34_add_66848_comb;
  wire [31:0] p34_add_66869_comb;
  wire [31:0] p34_add_66904_comb;
  wire [31:0] p34_add_66905_comb;
  wire [31:0] p34_add_66809_comb;
  wire [31:0] p34_add_66815_comb;
  wire [31:0] p34_add_66849_comb;
  wire [31:0] p34_add_66893_comb;
  wire [31:0] p34_add_66906_comb;
  assign p34_and_66850_comb = p33_add_66735 & p33_add_66633;
  assign p34_add_66807_comb = (p33_add_66707 & p33_add_66608 ^ ~(p33_add_66707 | ~p33_add_66509)) + {p33_add_66707[5:0] ^ p33_add_66707[10:5] ^ p33_add_66707[24:19], p33_add_66707[31:27] ^ p33_add_66707[4:0] ^ p33_add_66707[18:14], p33_add_66707[26:13] ^ p33_add_66707[31:18] ^ p33_add_66707[13:0], p33_add_66707[12:6] ^ p33_add_66707[17:11] ^ p33_add_66707[31:25]};
  assign p34_add_66812_comb = p33_add_65186[31:2] + 30'h134b_1b7f;
  assign p34_add_66808_comb = p34_add_66807_comb + p33_add_66713;
  assign p34_add_66847_comb = p33_add_64613 + {p33_add_64256[6:4] ^ p33_add_64256[17:15], p33_add_64256[3:0] ^ p33_add_64256[14:11] ^ p33_add_64256[31:28], p33_add_64256[31:21] ^ p33_add_64256[10:0] ^ p33_add_64256[27:17], p33_add_64256[20:7] ^ p33_add_64256[31:18] ^ p33_add_64256[16:3]};
  assign p34_add_66848_comb = {p33_add_65186[16:7] ^ p33_add_65186[18:9], p33_add_65186[6:0] ^ p33_add_65186[8:2] ^ p33_add_65186[31:25], p33_add_65186[31:30] ^ p33_add_65186[1:0] ^ p33_add_65186[24:23], p33_add_65186[29:17] ^ p33_add_65186[31:19] ^ p33_add_65186[22:10]} + p33_add_63929;
  assign p34_add_66869_comb = (p34_and_66850_comb ^ p33_add_66735 & p33_add_66534 ^ p33_and_66714) + p33_add_66706;
  assign p34_add_66904_comb = p33_add_64631 + {p33_add_63999[6:4] ^ p33_add_63999[17:15], p33_add_63999[3:0] ^ p33_add_63999[14:11] ^ p33_add_63999[31:28], p33_add_63999[31:21] ^ p33_add_63999[10:0] ^ p33_add_63999[27:17], p33_add_63999[20:7] ^ p33_add_63999[31:18] ^ p33_add_63999[16:3]};
  assign p34_add_66905_comb = {p33_add_65326[16:7] ^ p33_add_65326[18:9], p33_add_65326[6:0] ^ p33_add_65326[8:2] ^ p33_add_65326[31:25], p33_add_65326[31:30] ^ p33_add_65326[1:0] ^ p33_add_65326[24:23], p33_add_65326[29:17] ^ p33_add_65326[31:19] ^ p33_add_65326[22:10]} + p33_add_64256;
  assign p34_add_66809_comb = p34_add_66808_comb + p33_add_66534;
  assign p34_add_66815_comb = {p34_add_66812_comb, p33_add_65186[1:0]} + p33_add_66509;
  assign p34_add_66849_comb = p34_add_66847_comb + p34_add_66848_comb;
  assign p34_add_66893_comb = p34_add_66869_comb + {p33_add_66735[1:0] ^ p33_add_66735[12:11] ^ p33_add_66735[21:20], p33_add_66735[31:21] ^ p33_add_66735[10:0] ^ p33_add_66735[19:9], p33_add_66735[20:12] ^ p33_add_66735[31:23] ^ p33_add_66735[8:0], p33_add_66735[11:2] ^ p33_add_66735[22:13] ^ p33_add_66735[31:22]};
  assign p34_add_66906_comb = p34_add_66904_comb + p34_add_66905_comb;

  // Registers for pipe stage 34:
  reg [31:0] p34_add_63999;
  reg [31:0] p34_add_64275;
  reg [31:0] p34_add_64292;
  reg [31:0] p34_add_64444;
  reg [31:0] p34_add_64445;
  reg [31:0] p34_add_64595;
  reg [31:0] p34_add_64480;
  reg [31:0] p34_add_64613;
  reg [31:0] p34_add_64631;
  reg [31:0] p34_add_64766;
  reg [31:0] p34_add_66608;
  reg [31:0] p34_add_64904;
  reg [31:0] p34_add_66707;
  reg [31:0] p34_add_65045;
  reg [31:0] p34_add_66808;
  reg [31:0] p34_add_66809;
  reg [31:0] p34_add_65186;
  reg [31:0] p34_add_66815;
  reg [31:0] p34_add_66633;
  reg [31:0] p34_add_65326;
  reg [31:0] p34_add_66735;
  reg [31:0] p34_add_66849;
  reg [31:0] p34_and_66850;
  reg [31:0] p34_add_66893;
  reg [31:0] p34_add_66906;
  always_ff @ (posedge clk) begin
    p34_add_63999 <= p33_add_63999;
    p34_add_64275 <= p33_add_64275;
    p34_add_64292 <= p33_add_64292;
    p34_add_64444 <= p33_add_64444;
    p34_add_64445 <= p33_add_64445;
    p34_add_64595 <= p33_add_64595;
    p34_add_64480 <= p33_add_64480;
    p34_add_64613 <= p33_add_64613;
    p34_add_64631 <= p33_add_64631;
    p34_add_64766 <= p33_add_64766;
    p34_add_66608 <= p33_add_66608;
    p34_add_64904 <= p33_add_64904;
    p34_add_66707 <= p33_add_66707;
    p34_add_65045 <= p33_add_65045;
    p34_add_66808 <= p34_add_66808_comb;
    p34_add_66809 <= p34_add_66809_comb;
    p34_add_65186 <= p33_add_65186;
    p34_add_66815 <= p34_add_66815_comb;
    p34_add_66633 <= p33_add_66633;
    p34_add_65326 <= p33_add_65326;
    p34_add_66735 <= p33_add_66735;
    p34_add_66849 <= p34_add_66849_comb;
    p34_and_66850 <= p34_and_66850_comb;
    p34_add_66893 <= p34_add_66893_comb;
    p34_add_66906 <= p34_add_66906_comb;
  end

  // ===== Pipe stage 35:
  wire [1:0] p35_bit_slice_66984_comb;
  wire [31:0] p35_add_67038_comb;
  wire [31:0] p35_add_67039_comb;
  wire [31:0] p35_add_67040_comb;
  wire [31:0] p35_and_66985_comb;
  wire [31:0] p35_add_66978_comb;
  wire [31:0] p35_add_66979_comb;
  wire [31:0] p35_add_66982_comb;
  wire [31:0] p35_add_67033_comb;
  wire [31:0] p35_add_67073_comb;
  wire [31:0] p35_add_67074_comb;
  wire [31:0] p35_add_66980_comb;
  wire [31:0] p35_add_66983_comb;
  wire [31:0] p35_add_67037_comb;
  wire [31:0] p35_add_67075_comb;
  wire [31:0] p35_add_67092_comb;
  assign p35_bit_slice_66984_comb = p34_add_66849[1:0];
  assign p35_add_67038_comb = p34_add_64766 + {p34_add_64275[6:4] ^ p34_add_64275[17:15], p34_add_64275[3:0] ^ p34_add_64275[14:11] ^ p34_add_64275[31:28], p34_add_64275[31:21] ^ p34_add_64275[10:0] ^ p34_add_64275[27:17], p34_add_64275[20:7] ^ p34_add_64275[31:18] ^ p34_add_64275[16:3]};
  assign p35_add_67039_comb = {p34_add_66849[16:7] ^ p34_add_66849[18:9], p34_add_66849[6:0] ^ p34_add_66849[8:2] ^ p34_add_66849[31:25], p34_add_66849[31:30] ^ p35_bit_slice_66984_comb ^ p34_add_66849[24:23], p34_add_66849[29:17] ^ p34_add_66849[31:19] ^ p34_add_66849[22:10]} + p34_add_63999;
  assign p35_add_67040_comb = p35_add_67038_comb + p35_add_67039_comb;
  assign p35_and_66985_comb = p34_add_66893 & p34_add_66735;
  assign p35_add_66978_comb = (p34_add_66809 & p34_add_66707 ^ ~(p34_add_66809 | ~p34_add_66608)) + {p34_add_66809[5:0] ^ p34_add_66809[10:5] ^ p34_add_66809[24:19], p34_add_66809[31:27] ^ p34_add_66809[4:0] ^ p34_add_66809[18:14], p34_add_66809[26:13] ^ p34_add_66809[31:18] ^ p34_add_66809[13:0], p34_add_66809[12:6] ^ p34_add_66809[17:11] ^ p34_add_66809[31:25]};
  assign p35_add_66979_comb = p35_add_66978_comb + p34_add_66815;
  assign p35_add_66982_comb = p34_add_65326 + 32'h5338_0d13;
  assign p35_add_67033_comb = (p35_and_66985_comb ^ p34_add_66893 & p34_add_66633 ^ p34_and_66850) + p34_add_66808;
  assign p35_add_67073_comb = p34_add_64904 + {p34_add_64292[6:4] ^ p34_add_64292[17:15], p34_add_64292[3:0] ^ p34_add_64292[14:11] ^ p34_add_64292[31:28], p34_add_64292[31:21] ^ p34_add_64292[10:0] ^ p34_add_64292[27:17], p34_add_64292[20:7] ^ p34_add_64292[31:18] ^ p34_add_64292[16:3]};
  assign p35_add_67074_comb = {p34_add_66906[16:7] ^ p34_add_66906[18:9], p34_add_66906[6:0] ^ p34_add_66906[8:2] ^ p34_add_66906[31:25], p34_add_66906[31:30] ^ p34_add_66906[1:0] ^ p34_add_66906[24:23], p34_add_66906[29:17] ^ p34_add_66906[31:19] ^ p34_add_66906[22:10]} + p34_add_64275;
  assign p35_add_66980_comb = p35_add_66979_comb + p34_add_66633;
  assign p35_add_66983_comb = p34_add_66608 + p35_add_66982_comb;
  assign p35_add_67037_comb = p35_add_67033_comb + {p34_add_66893[1:0] ^ p34_add_66893[12:11] ^ p34_add_66893[21:20], p34_add_66893[31:21] ^ p34_add_66893[10:0] ^ p34_add_66893[19:9], p34_add_66893[20:12] ^ p34_add_66893[31:23] ^ p34_add_66893[8:0], p34_add_66893[11:2] ^ p34_add_66893[22:13] ^ p34_add_66893[31:22]};
  assign p35_add_67075_comb = p35_add_67073_comb + p35_add_67074_comb;
  assign p35_add_67092_comb = {p35_add_67040_comb[16:7] ^ p35_add_67040_comb[18:9], p35_add_67040_comb[6:0] ^ p35_add_67040_comb[8:2] ^ p35_add_67040_comb[31:25], p35_add_67040_comb[31:30] ^ p35_add_67040_comb[1:0] ^ p35_add_67040_comb[24:23], p35_add_67040_comb[29:17] ^ p35_add_67040_comb[31:19] ^ p35_add_67040_comb[22:10]} + p34_add_64292;

  // Registers for pipe stage 35:
  reg [31:0] p35_add_64444;
  reg [31:0] p35_add_64445;
  reg [31:0] p35_add_64595;
  reg [31:0] p35_add_64480;
  reg [31:0] p35_add_64613;
  reg [31:0] p35_add_64631;
  reg [31:0] p35_add_64766;
  reg [31:0] p35_add_64904;
  reg [31:0] p35_add_66707;
  reg [31:0] p35_add_65045;
  reg [31:0] p35_add_66809;
  reg [31:0] p35_add_65186;
  reg [31:0] p35_add_66979;
  reg [31:0] p35_add_66980;
  reg [31:0] p35_add_65326;
  reg [31:0] p35_add_66983;
  reg [31:0] p35_add_66735;
  reg [31:0] p35_add_66849;
  reg [1:0] p35_bit_slice_66984;
  reg [31:0] p35_add_66893;
  reg [31:0] p35_add_66906;
  reg [31:0] p35_and_66985;
  reg [31:0] p35_add_67037;
  reg [31:0] p35_add_67040;
  reg [31:0] p35_add_67075;
  reg [31:0] p35_add_67092;
  always_ff @ (posedge clk) begin
    p35_add_64444 <= p34_add_64444;
    p35_add_64445 <= p34_add_64445;
    p35_add_64595 <= p34_add_64595;
    p35_add_64480 <= p34_add_64480;
    p35_add_64613 <= p34_add_64613;
    p35_add_64631 <= p34_add_64631;
    p35_add_64766 <= p34_add_64766;
    p35_add_64904 <= p34_add_64904;
    p35_add_66707 <= p34_add_66707;
    p35_add_65045 <= p34_add_65045;
    p35_add_66809 <= p34_add_66809;
    p35_add_65186 <= p34_add_65186;
    p35_add_66979 <= p35_add_66979_comb;
    p35_add_66980 <= p35_add_66980_comb;
    p35_add_65326 <= p34_add_65326;
    p35_add_66983 <= p35_add_66983_comb;
    p35_add_66735 <= p34_add_66735;
    p35_add_66849 <= p34_add_66849;
    p35_bit_slice_66984 <= p35_bit_slice_66984_comb;
    p35_add_66893 <= p34_add_66893;
    p35_add_66906 <= p34_add_66906;
    p35_and_66985 <= p35_and_66985_comb;
    p35_add_67037 <= p35_add_67037_comb;
    p35_add_67040 <= p35_add_67040_comb;
    p35_add_67075 <= p35_add_67075_comb;
    p35_add_67092 <= p35_add_67092_comb;
  end

  // ===== Pipe stage 36:
  wire [31:0] p36_add_67212_comb;
  wire [31:0] p36_add_67213_comb;
  wire [31:0] p36_and_67174_comb;
  wire [31:0] p36_add_67166_comb;
  wire [29:0] p36_add_67171_comb;
  wire [31:0] p36_add_67167_comb;
  wire [31:0] p36_add_67193_comb;
  wire [31:0] p36_add_67246_comb;
  wire [31:0] p36_add_67247_comb;
  wire [31:0] p36_add_67168_comb;
  wire [31:0] p36_add_67173_comb;
  wire [31:0] p36_add_67195_comb;
  wire [31:0] p36_add_67248_comb;
  wire [31:0] p36_add_67265_comb;
  assign p36_add_67212_comb = p35_add_65045 + {p35_add_64444[6:4] ^ p35_add_64444[17:15], p35_add_64444[3:0] ^ p35_add_64444[14:11] ^ p35_add_64444[31:28], p35_add_64444[31:21] ^ p35_add_64444[10:0] ^ p35_add_64444[27:17], p35_add_64444[20:7] ^ p35_add_64444[31:18] ^ p35_add_64444[16:3]};
  assign p36_add_67213_comb = p36_add_67212_comb + p35_add_67092;
  assign p36_and_67174_comb = p35_add_67037 & p35_add_66893;
  assign p36_add_67166_comb = {p35_add_66980[5:0] ^ p35_add_66980[10:5] ^ p35_add_66980[24:19], p35_add_66980[31:27] ^ p35_add_66980[4:0] ^ p35_add_66980[18:14], p35_add_66980[26:13] ^ p35_add_66980[31:18] ^ p35_add_66980[13:0], p35_add_66980[12:6] ^ p35_add_66980[17:11] ^ p35_add_66980[31:25]} + (p35_add_66980 & p35_add_66809 ^ ~(p35_add_66980 | ~p35_add_66707));
  assign p36_add_67171_comb = p35_add_66849[31:2] + 30'h1942_9cd5;
  assign p36_add_67167_comb = p36_add_67166_comb + p35_add_66983;
  assign p36_add_67193_comb = (p36_and_67174_comb ^ p35_add_67037 & p35_add_66735 ^ p35_and_66985) + p35_add_66979;
  assign p36_add_67246_comb = p35_add_65186 + {p35_add_64445[6:4] ^ p35_add_64445[17:15], p35_add_64445[3:0] ^ p35_add_64445[14:11] ^ p35_add_64445[31:28], p35_add_64445[31:21] ^ p35_add_64445[10:0] ^ p35_add_64445[27:17], p35_add_64445[20:7] ^ p35_add_64445[31:18] ^ p35_add_64445[16:3]};
  assign p36_add_67247_comb = {p35_add_67075[16:7] ^ p35_add_67075[18:9], p35_add_67075[6:0] ^ p35_add_67075[8:2] ^ p35_add_67075[31:25], p35_add_67075[31:30] ^ p35_add_67075[1:0] ^ p35_add_67075[24:23], p35_add_67075[29:17] ^ p35_add_67075[31:19] ^ p35_add_67075[22:10]} + p35_add_64444;
  assign p36_add_67168_comb = p36_add_67167_comb + p35_add_66735;
  assign p36_add_67173_comb = {p36_add_67171_comb, p35_bit_slice_66984} + p35_add_66707;
  assign p36_add_67195_comb = p36_add_67193_comb + {p35_add_67037[1:0] ^ p35_add_67037[12:11] ^ p35_add_67037[21:20], p35_add_67037[31:21] ^ p35_add_67037[10:0] ^ p35_add_67037[19:9], p35_add_67037[20:12] ^ p35_add_67037[31:23] ^ p35_add_67037[8:0], p35_add_67037[11:2] ^ p35_add_67037[22:13] ^ p35_add_67037[31:22]};
  assign p36_add_67248_comb = p36_add_67246_comb + p36_add_67247_comb;
  assign p36_add_67265_comb = {p36_add_67213_comb[16:7] ^ p36_add_67213_comb[18:9], p36_add_67213_comb[6:0] ^ p36_add_67213_comb[8:2] ^ p36_add_67213_comb[31:25], p36_add_67213_comb[31:30] ^ p36_add_67213_comb[1:0] ^ p36_add_67213_comb[24:23], p36_add_67213_comb[29:17] ^ p36_add_67213_comb[31:19] ^ p36_add_67213_comb[22:10]} + p35_add_64445;

  // Registers for pipe stage 36:
  reg [31:0] p36_add_64595;
  reg [31:0] p36_add_64480;
  reg [31:0] p36_add_64613;
  reg [31:0] p36_add_64631;
  reg [31:0] p36_add_64766;
  reg [31:0] p36_add_64904;
  reg [31:0] p36_add_65045;
  reg [31:0] p36_add_66809;
  reg [31:0] p36_add_65186;
  reg [31:0] p36_add_66980;
  reg [31:0] p36_add_65326;
  reg [31:0] p36_add_67167;
  reg [31:0] p36_add_67168;
  reg [31:0] p36_add_66849;
  reg [31:0] p36_add_67173;
  reg [31:0] p36_add_66893;
  reg [31:0] p36_add_66906;
  reg [31:0] p36_add_67037;
  reg [31:0] p36_add_67040;
  reg [31:0] p36_and_67174;
  reg [31:0] p36_add_67195;
  reg [31:0] p36_add_67075;
  reg [31:0] p36_add_67213;
  reg [31:0] p36_add_67248;
  reg [31:0] p36_add_67265;
  always_ff @ (posedge clk) begin
    p36_add_64595 <= p35_add_64595;
    p36_add_64480 <= p35_add_64480;
    p36_add_64613 <= p35_add_64613;
    p36_add_64631 <= p35_add_64631;
    p36_add_64766 <= p35_add_64766;
    p36_add_64904 <= p35_add_64904;
    p36_add_65045 <= p35_add_65045;
    p36_add_66809 <= p35_add_66809;
    p36_add_65186 <= p35_add_65186;
    p36_add_66980 <= p35_add_66980;
    p36_add_65326 <= p35_add_65326;
    p36_add_67167 <= p36_add_67167_comb;
    p36_add_67168 <= p36_add_67168_comb;
    p36_add_66849 <= p35_add_66849;
    p36_add_67173 <= p36_add_67173_comb;
    p36_add_66893 <= p35_add_66893;
    p36_add_66906 <= p35_add_66906;
    p36_add_67037 <= p35_add_67037;
    p36_add_67040 <= p35_add_67040;
    p36_and_67174 <= p36_and_67174_comb;
    p36_add_67195 <= p36_add_67195_comb;
    p36_add_67075 <= p35_add_67075;
    p36_add_67213 <= p36_add_67213_comb;
    p36_add_67248 <= p36_add_67248_comb;
    p36_add_67265 <= p36_add_67265_comb;
  end

  // ===== Pipe stage 37:
  wire [31:0] p37_add_67381_comb;
  wire [31:0] p37_add_67382_comb;
  wire [31:0] p37_and_67343_comb;
  wire [31:0] p37_add_67337_comb;
  wire [31:0] p37_add_67338_comb;
  wire [31:0] p37_add_67341_comb;
  wire [31:0] p37_add_67362_comb;
  wire [31:0] p37_add_67415_comb;
  wire [31:0] p37_add_67416_comb;
  wire [31:0] p37_add_67339_comb;
  wire [31:0] p37_add_67342_comb;
  wire [31:0] p37_add_67364_comb;
  wire [31:0] p37_add_67417_comb;
  wire [31:0] p37_add_67434_comb;
  assign p37_add_67381_comb = p36_add_65326 + {p36_add_64595[6:4] ^ p36_add_64595[17:15], p36_add_64595[3:0] ^ p36_add_64595[14:11] ^ p36_add_64595[31:28], p36_add_64595[31:21] ^ p36_add_64595[10:0] ^ p36_add_64595[27:17], p36_add_64595[20:7] ^ p36_add_64595[31:18] ^ p36_add_64595[16:3]};
  assign p37_add_67382_comb = p37_add_67381_comb + p36_add_67265;
  assign p37_and_67343_comb = p36_add_67195 & p36_add_67037;
  assign p37_add_67337_comb = (p36_add_67168 & p36_add_66980 ^ ~(p36_add_67168 | ~p36_add_66809)) + {p36_add_67168[5:0] ^ p36_add_67168[10:5] ^ p36_add_67168[24:19], p36_add_67168[31:27] ^ p36_add_67168[4:0] ^ p36_add_67168[18:14], p36_add_67168[26:13] ^ p36_add_67168[31:18] ^ p36_add_67168[13:0], p36_add_67168[12:6] ^ p36_add_67168[17:11] ^ p36_add_67168[31:25]};
  assign p37_add_67338_comb = p37_add_67337_comb + p36_add_67173;
  assign p37_add_67341_comb = p36_add_66906 + 32'h766a_0abb;
  assign p37_add_67362_comb = (p37_and_67343_comb ^ p36_add_67195 & p36_add_66893 ^ p36_and_67174) + p36_add_67167;
  assign p37_add_67415_comb = p36_add_66849 + {p36_add_64480[6:4] ^ p36_add_64480[17:15], p36_add_64480[3:0] ^ p36_add_64480[14:11] ^ p36_add_64480[31:28], p36_add_64480[31:21] ^ p36_add_64480[10:0] ^ p36_add_64480[27:17], p36_add_64480[20:7] ^ p36_add_64480[31:18] ^ p36_add_64480[16:3]};
  assign p37_add_67416_comb = {p36_add_67248[16:7] ^ p36_add_67248[18:9], p36_add_67248[6:0] ^ p36_add_67248[8:2] ^ p36_add_67248[31:25], p36_add_67248[31:30] ^ p36_add_67248[1:0] ^ p36_add_67248[24:23], p36_add_67248[29:17] ^ p36_add_67248[31:19] ^ p36_add_67248[22:10]} + p36_add_64595;
  assign p37_add_67339_comb = p37_add_67338_comb + p36_add_66893;
  assign p37_add_67342_comb = p36_add_66809 + p37_add_67341_comb;
  assign p37_add_67364_comb = p37_add_67362_comb + {p36_add_67195[1:0] ^ p36_add_67195[12:11] ^ p36_add_67195[21:20], p36_add_67195[31:21] ^ p36_add_67195[10:0] ^ p36_add_67195[19:9], p36_add_67195[20:12] ^ p36_add_67195[31:23] ^ p36_add_67195[8:0], p36_add_67195[11:2] ^ p36_add_67195[22:13] ^ p36_add_67195[31:22]};
  assign p37_add_67417_comb = p37_add_67415_comb + p37_add_67416_comb;
  assign p37_add_67434_comb = {p37_add_67382_comb[16:7] ^ p37_add_67382_comb[18:9], p37_add_67382_comb[6:0] ^ p37_add_67382_comb[8:2] ^ p37_add_67382_comb[31:25], p37_add_67382_comb[31:30] ^ p37_add_67382_comb[1:0] ^ p37_add_67382_comb[24:23], p37_add_67382_comb[29:17] ^ p37_add_67382_comb[31:19] ^ p37_add_67382_comb[22:10]} + p36_add_64480;

  // Registers for pipe stage 37:
  reg [31:0] p37_add_64613;
  reg [31:0] p37_add_64631;
  reg [31:0] p37_add_64766;
  reg [31:0] p37_add_64904;
  reg [31:0] p37_add_65045;
  reg [31:0] p37_add_65186;
  reg [31:0] p37_add_66980;
  reg [31:0] p37_add_65326;
  reg [31:0] p37_add_67168;
  reg [31:0] p37_add_66849;
  reg [31:0] p37_add_67338;
  reg [31:0] p37_add_67339;
  reg [31:0] p37_add_66906;
  reg [31:0] p37_add_67342;
  reg [31:0] p37_add_67037;
  reg [31:0] p37_add_67040;
  reg [31:0] p37_add_67195;
  reg [31:0] p37_add_67075;
  reg [31:0] p37_and_67343;
  reg [31:0] p37_add_67364;
  reg [31:0] p37_add_67213;
  reg [31:0] p37_add_67248;
  reg [31:0] p37_add_67382;
  reg [31:0] p37_add_67417;
  reg [31:0] p37_add_67434;
  always_ff @ (posedge clk) begin
    p37_add_64613 <= p36_add_64613;
    p37_add_64631 <= p36_add_64631;
    p37_add_64766 <= p36_add_64766;
    p37_add_64904 <= p36_add_64904;
    p37_add_65045 <= p36_add_65045;
    p37_add_65186 <= p36_add_65186;
    p37_add_66980 <= p36_add_66980;
    p37_add_65326 <= p36_add_65326;
    p37_add_67168 <= p36_add_67168;
    p37_add_66849 <= p36_add_66849;
    p37_add_67338 <= p37_add_67338_comb;
    p37_add_67339 <= p37_add_67339_comb;
    p37_add_66906 <= p36_add_66906;
    p37_add_67342 <= p37_add_67342_comb;
    p37_add_67037 <= p36_add_67037;
    p37_add_67040 <= p36_add_67040;
    p37_add_67195 <= p36_add_67195;
    p37_add_67075 <= p36_add_67075;
    p37_and_67343 <= p37_and_67343_comb;
    p37_add_67364 <= p37_add_67364_comb;
    p37_add_67213 <= p36_add_67213;
    p37_add_67248 <= p36_add_67248;
    p37_add_67382 <= p37_add_67382_comb;
    p37_add_67417 <= p37_add_67417_comb;
    p37_add_67434 <= p37_add_67434_comb;
  end

  // ===== Pipe stage 38:
  wire [31:0] p38_add_67553_comb;
  wire [31:0] p38_add_67554_comb;
  wire [31:0] p38_and_67515_comb;
  wire [31:0] p38_add_67506_comb;
  wire [30:0] p38_add_67511_comb;
  wire [31:0] p38_add_67507_comb;
  wire [31:0] p38_add_67534_comb;
  wire [31:0] p38_add_67587_comb;
  wire [31:0] p38_add_67588_comb;
  wire [31:0] p38_add_67508_comb;
  wire [31:0] p38_add_67514_comb;
  wire [31:0] p38_add_67536_comb;
  wire [31:0] p38_add_67589_comb;
  wire [31:0] p38_add_67606_comb;
  assign p38_add_67553_comb = p37_add_66906 + {p37_add_64613[6:4] ^ p37_add_64613[17:15], p37_add_64613[3:0] ^ p37_add_64613[14:11] ^ p37_add_64613[31:28], p37_add_64613[31:21] ^ p37_add_64613[10:0] ^ p37_add_64613[27:17], p37_add_64613[20:7] ^ p37_add_64613[31:18] ^ p37_add_64613[16:3]};
  assign p38_add_67554_comb = p38_add_67553_comb + p37_add_67434;
  assign p38_and_67515_comb = p37_add_67364 & p37_add_67195;
  assign p38_add_67506_comb = {p37_add_67339[5:0] ^ p37_add_67339[10:5] ^ p37_add_67339[24:19], p37_add_67339[31:27] ^ p37_add_67339[4:0] ^ p37_add_67339[18:14], p37_add_67339[26:13] ^ p37_add_67339[31:18] ^ p37_add_67339[13:0], p37_add_67339[12:6] ^ p37_add_67339[17:11] ^ p37_add_67339[31:25]} + (p37_add_67339 & p37_add_67168 ^ ~(p37_add_67339 | ~p37_add_66980));
  assign p38_add_67511_comb = p37_add_67040[31:1] + 31'h40e1_6497;
  assign p38_add_67507_comb = p38_add_67506_comb + p37_add_67342;
  assign p38_add_67534_comb = (p38_and_67515_comb ^ p37_add_67364 & p37_add_67037 ^ p37_and_67343) + p37_add_67338;
  assign p38_add_67587_comb = p37_add_67040 + {p37_add_64631[6:4] ^ p37_add_64631[17:15], p37_add_64631[3:0] ^ p37_add_64631[14:11] ^ p37_add_64631[31:28], p37_add_64631[31:21] ^ p37_add_64631[10:0] ^ p37_add_64631[27:17], p37_add_64631[20:7] ^ p37_add_64631[31:18] ^ p37_add_64631[16:3]};
  assign p38_add_67588_comb = {p37_add_67417[16:7] ^ p37_add_67417[18:9], p37_add_67417[6:0] ^ p37_add_67417[8:2] ^ p37_add_67417[31:25], p37_add_67417[31:30] ^ p37_add_67417[1:0] ^ p37_add_67417[24:23], p37_add_67417[29:17] ^ p37_add_67417[31:19] ^ p37_add_67417[22:10]} + p37_add_64613;
  assign p38_add_67508_comb = p38_add_67507_comb + p37_add_67037;
  assign p38_add_67514_comb = {p38_add_67511_comb, p37_add_67040[0]} + p37_add_66980;
  assign p38_add_67536_comb = p38_add_67534_comb + {p37_add_67364[1:0] ^ p37_add_67364[12:11] ^ p37_add_67364[21:20], p37_add_67364[31:21] ^ p37_add_67364[10:0] ^ p37_add_67364[19:9], p37_add_67364[20:12] ^ p37_add_67364[31:23] ^ p37_add_67364[8:0], p37_add_67364[11:2] ^ p37_add_67364[22:13] ^ p37_add_67364[31:22]};
  assign p38_add_67589_comb = p38_add_67587_comb + p38_add_67588_comb;
  assign p38_add_67606_comb = {p38_add_67554_comb[16:7] ^ p38_add_67554_comb[18:9], p38_add_67554_comb[6:0] ^ p38_add_67554_comb[8:2] ^ p38_add_67554_comb[31:25], p38_add_67554_comb[31:30] ^ p38_add_67554_comb[1:0] ^ p38_add_67554_comb[24:23], p38_add_67554_comb[29:17] ^ p38_add_67554_comb[31:19] ^ p38_add_67554_comb[22:10]} + p37_add_64631;

  // Registers for pipe stage 38:
  reg [31:0] p38_add_64766;
  reg [31:0] p38_add_64904;
  reg [31:0] p38_add_65045;
  reg [31:0] p38_add_65186;
  reg [31:0] p38_add_65326;
  reg [31:0] p38_add_67168;
  reg [31:0] p38_add_66849;
  reg [31:0] p38_add_67339;
  reg [31:0] p38_add_66906;
  reg [31:0] p38_add_67507;
  reg [31:0] p38_add_67508;
  reg [31:0] p38_add_67040;
  reg [31:0] p38_add_67514;
  reg [31:0] p38_add_67195;
  reg [31:0] p38_add_67075;
  reg [31:0] p38_add_67364;
  reg [31:0] p38_add_67213;
  reg [31:0] p38_and_67515;
  reg [31:0] p38_add_67536;
  reg [31:0] p38_add_67248;
  reg [31:0] p38_add_67382;
  reg [31:0] p38_add_67417;
  reg [31:0] p38_add_67554;
  reg [31:0] p38_add_67589;
  reg [31:0] p38_add_67606;
  always_ff @ (posedge clk) begin
    p38_add_64766 <= p37_add_64766;
    p38_add_64904 <= p37_add_64904;
    p38_add_65045 <= p37_add_65045;
    p38_add_65186 <= p37_add_65186;
    p38_add_65326 <= p37_add_65326;
    p38_add_67168 <= p37_add_67168;
    p38_add_66849 <= p37_add_66849;
    p38_add_67339 <= p37_add_67339;
    p38_add_66906 <= p37_add_66906;
    p38_add_67507 <= p38_add_67507_comb;
    p38_add_67508 <= p38_add_67508_comb;
    p38_add_67040 <= p37_add_67040;
    p38_add_67514 <= p38_add_67514_comb;
    p38_add_67195 <= p37_add_67195;
    p38_add_67075 <= p37_add_67075;
    p38_add_67364 <= p37_add_67364;
    p38_add_67213 <= p37_add_67213;
    p38_and_67515 <= p38_and_67515_comb;
    p38_add_67536 <= p38_add_67536_comb;
    p38_add_67248 <= p37_add_67248;
    p38_add_67382 <= p37_add_67382;
    p38_add_67417 <= p37_add_67417;
    p38_add_67554 <= p38_add_67554_comb;
    p38_add_67589 <= p38_add_67589_comb;
    p38_add_67606 <= p38_add_67606_comb;
  end

  // ===== Pipe stage 39:
  wire [31:0] p39_add_67723_comb;
  wire [1:0] p39_bit_slice_67706_comb;
  wire [31:0] p39_add_67724_comb;
  wire [31:0] p39_and_67684_comb;
  wire [31:0] p39_add_67678_comb;
  wire [31:0] p39_add_67679_comb;
  wire [31:0] p39_add_67682_comb;
  wire [31:0] p39_add_67703_comb;
  wire [31:0] p39_add_67756_comb;
  wire [31:0] p39_add_67757_comb;
  wire [31:0] p39_add_67680_comb;
  wire [31:0] p39_add_67683_comb;
  wire [31:0] p39_add_67705_comb;
  wire [31:0] p39_add_67758_comb;
  wire [31:0] p39_add_67775_comb;
  assign p39_add_67723_comb = p38_add_67075 + {p38_add_64766[6:4] ^ p38_add_64766[17:15], p38_add_64766[3:0] ^ p38_add_64766[14:11] ^ p38_add_64766[31:28], p38_add_64766[31:21] ^ p38_add_64766[10:0] ^ p38_add_64766[27:17], p38_add_64766[20:7] ^ p38_add_64766[31:18] ^ p38_add_64766[16:3]};
  assign p39_bit_slice_67706_comb = p38_add_67589[1:0];
  assign p39_add_67724_comb = p39_add_67723_comb + p38_add_67606;
  assign p39_and_67684_comb = p38_add_67536 & p38_add_67364;
  assign p39_add_67678_comb = (p38_add_67508 & p38_add_67339 ^ ~(p38_add_67508 | ~p38_add_67168)) + {p38_add_67508[5:0] ^ p38_add_67508[10:5] ^ p38_add_67508[24:19], p38_add_67508[31:27] ^ p38_add_67508[4:0] ^ p38_add_67508[18:14], p38_add_67508[26:13] ^ p38_add_67508[31:18] ^ p38_add_67508[13:0], p38_add_67508[12:6] ^ p38_add_67508[17:11] ^ p38_add_67508[31:25]};
  assign p39_add_67679_comb = p39_add_67678_comb + p38_add_67514;
  assign p39_add_67682_comb = p38_add_67075 + 32'h9272_2c85;
  assign p39_add_67703_comb = (p39_and_67684_comb ^ p38_add_67536 & p38_add_67195 ^ p38_and_67515) + p38_add_67507;
  assign p39_add_67756_comb = p38_add_67213 + {p38_add_64904[6:4] ^ p38_add_64904[17:15], p38_add_64904[3:0] ^ p38_add_64904[14:11] ^ p38_add_64904[31:28], p38_add_64904[31:21] ^ p38_add_64904[10:0] ^ p38_add_64904[27:17], p38_add_64904[20:7] ^ p38_add_64904[31:18] ^ p38_add_64904[16:3]};
  assign p39_add_67757_comb = {p38_add_67589[16:7] ^ p38_add_67589[18:9], p38_add_67589[6:0] ^ p38_add_67589[8:2] ^ p38_add_67589[31:25], p38_add_67589[31:30] ^ p39_bit_slice_67706_comb ^ p38_add_67589[24:23], p38_add_67589[29:17] ^ p38_add_67589[31:19] ^ p38_add_67589[22:10]} + p38_add_64766;
  assign p39_add_67680_comb = p39_add_67679_comb + p38_add_67195;
  assign p39_add_67683_comb = p38_add_67168 + p39_add_67682_comb;
  assign p39_add_67705_comb = p39_add_67703_comb + {p38_add_67536[1:0] ^ p38_add_67536[12:11] ^ p38_add_67536[21:20], p38_add_67536[31:21] ^ p38_add_67536[10:0] ^ p38_add_67536[19:9], p38_add_67536[20:12] ^ p38_add_67536[31:23] ^ p38_add_67536[8:0], p38_add_67536[11:2] ^ p38_add_67536[22:13] ^ p38_add_67536[31:22]};
  assign p39_add_67758_comb = p39_add_67756_comb + p39_add_67757_comb;
  assign p39_add_67775_comb = {p39_add_67724_comb[16:7] ^ p39_add_67724_comb[18:9], p39_add_67724_comb[6:0] ^ p39_add_67724_comb[8:2] ^ p39_add_67724_comb[31:25], p39_add_67724_comb[31:30] ^ p39_add_67724_comb[1:0] ^ p39_add_67724_comb[24:23], p39_add_67724_comb[29:17] ^ p39_add_67724_comb[31:19] ^ p39_add_67724_comb[22:10]} + p38_add_64904;

  // Registers for pipe stage 39:
  reg [31:0] p39_add_65045;
  reg [31:0] p39_add_65186;
  reg [31:0] p39_add_65326;
  reg [31:0] p39_add_66849;
  reg [31:0] p39_add_67339;
  reg [31:0] p39_add_66906;
  reg [31:0] p39_add_67508;
  reg [31:0] p39_add_67040;
  reg [31:0] p39_add_67679;
  reg [31:0] p39_add_67680;
  reg [31:0] p39_add_67075;
  reg [31:0] p39_add_67683;
  reg [31:0] p39_add_67364;
  reg [31:0] p39_add_67213;
  reg [31:0] p39_add_67536;
  reg [31:0] p39_add_67248;
  reg [31:0] p39_and_67684;
  reg [31:0] p39_add_67705;
  reg [31:0] p39_add_67382;
  reg [31:0] p39_add_67417;
  reg [31:0] p39_add_67554;
  reg [31:0] p39_add_67589;
  reg [1:0] p39_bit_slice_67706;
  reg [31:0] p39_add_67724;
  reg [31:0] p39_add_67758;
  reg [31:0] p39_add_67775;
  always_ff @ (posedge clk) begin
    p39_add_65045 <= p38_add_65045;
    p39_add_65186 <= p38_add_65186;
    p39_add_65326 <= p38_add_65326;
    p39_add_66849 <= p38_add_66849;
    p39_add_67339 <= p38_add_67339;
    p39_add_66906 <= p38_add_66906;
    p39_add_67508 <= p38_add_67508;
    p39_add_67040 <= p38_add_67040;
    p39_add_67679 <= p39_add_67679_comb;
    p39_add_67680 <= p39_add_67680_comb;
    p39_add_67075 <= p38_add_67075;
    p39_add_67683 <= p39_add_67683_comb;
    p39_add_67364 <= p38_add_67364;
    p39_add_67213 <= p38_add_67213;
    p39_add_67536 <= p38_add_67536;
    p39_add_67248 <= p38_add_67248;
    p39_and_67684 <= p39_and_67684_comb;
    p39_add_67705 <= p39_add_67705_comb;
    p39_add_67382 <= p38_add_67382;
    p39_add_67417 <= p38_add_67417;
    p39_add_67554 <= p38_add_67554;
    p39_add_67589 <= p38_add_67589;
    p39_bit_slice_67706 <= p39_bit_slice_67706_comb;
    p39_add_67724 <= p39_add_67724_comb;
    p39_add_67758 <= p39_add_67758_comb;
    p39_add_67775 <= p39_add_67775_comb;
  end

  // ===== Pipe stage 40:
  wire [31:0] p40_add_67893_comb;
  wire [31:0] p40_add_67894_comb;
  wire [31:0] p40_and_67855_comb;
  wire [31:0] p40_add_67849_comb;
  wire [31:0] p40_add_67850_comb;
  wire [31:0] p40_add_67853_comb;
  wire [31:0] p40_add_67874_comb;
  wire [31:0] p40_add_67927_comb;
  wire [31:0] p40_add_67928_comb;
  wire [31:0] p40_add_67851_comb;
  wire [31:0] p40_add_67854_comb;
  wire [31:0] p40_add_67876_comb;
  wire [31:0] p40_add_67929_comb;
  wire [31:0] p40_add_67946_comb;
  assign p40_add_67893_comb = p39_add_67248 + {p39_add_65045[6:4] ^ p39_add_65045[17:15], p39_add_65045[3:0] ^ p39_add_65045[14:11] ^ p39_add_65045[31:28], p39_add_65045[31:21] ^ p39_add_65045[10:0] ^ p39_add_65045[27:17], p39_add_65045[20:7] ^ p39_add_65045[31:18] ^ p39_add_65045[16:3]};
  assign p40_add_67894_comb = p40_add_67893_comb + p39_add_67775;
  assign p40_and_67855_comb = p39_add_67705 & p39_add_67536;
  assign p40_add_67849_comb = {p39_add_67680[5:0] ^ p39_add_67680[10:5] ^ p39_add_67680[24:19], p39_add_67680[31:27] ^ p39_add_67680[4:0] ^ p39_add_67680[18:14], p39_add_67680[26:13] ^ p39_add_67680[31:18] ^ p39_add_67680[13:0], p39_add_67680[12:6] ^ p39_add_67680[17:11] ^ p39_add_67680[31:25]} + (p39_add_67680 & p39_add_67508 ^ ~(p39_add_67680 | ~p39_add_67339));
  assign p40_add_67850_comb = p40_add_67849_comb + p39_add_67683;
  assign p40_add_67853_comb = p39_add_67213 + 32'ha2bf_e8a1;
  assign p40_add_67874_comb = (p40_and_67855_comb ^ p39_add_67705 & p39_add_67364 ^ p39_and_67684) + p39_add_67679;
  assign p40_add_67927_comb = p39_add_67382 + {p39_add_65186[6:4] ^ p39_add_65186[17:15], p39_add_65186[3:0] ^ p39_add_65186[14:11] ^ p39_add_65186[31:28], p39_add_65186[31:21] ^ p39_add_65186[10:0] ^ p39_add_65186[27:17], p39_add_65186[20:7] ^ p39_add_65186[31:18] ^ p39_add_65186[16:3]};
  assign p40_add_67928_comb = {p39_add_67758[16:7] ^ p39_add_67758[18:9], p39_add_67758[6:0] ^ p39_add_67758[8:2] ^ p39_add_67758[31:25], p39_add_67758[31:30] ^ p39_add_67758[1:0] ^ p39_add_67758[24:23], p39_add_67758[29:17] ^ p39_add_67758[31:19] ^ p39_add_67758[22:10]} + p39_add_65045;
  assign p40_add_67851_comb = p40_add_67850_comb + p39_add_67364;
  assign p40_add_67854_comb = p39_add_67339 + p40_add_67853_comb;
  assign p40_add_67876_comb = p40_add_67874_comb + {p39_add_67705[1:0] ^ p39_add_67705[12:11] ^ p39_add_67705[21:20], p39_add_67705[31:21] ^ p39_add_67705[10:0] ^ p39_add_67705[19:9], p39_add_67705[20:12] ^ p39_add_67705[31:23] ^ p39_add_67705[8:0], p39_add_67705[11:2] ^ p39_add_67705[22:13] ^ p39_add_67705[31:22]};
  assign p40_add_67929_comb = p40_add_67927_comb + p40_add_67928_comb;
  assign p40_add_67946_comb = {p40_add_67894_comb[16:7] ^ p40_add_67894_comb[18:9], p40_add_67894_comb[6:0] ^ p40_add_67894_comb[8:2] ^ p40_add_67894_comb[31:25], p40_add_67894_comb[31:30] ^ p40_add_67894_comb[1:0] ^ p40_add_67894_comb[24:23], p40_add_67894_comb[29:17] ^ p40_add_67894_comb[31:19] ^ p40_add_67894_comb[22:10]} + p39_add_65186;

  // Registers for pipe stage 40:
  reg [31:0] p40_add_65326;
  reg [31:0] p40_add_66849;
  reg [31:0] p40_add_66906;
  reg [31:0] p40_add_67508;
  reg [31:0] p40_add_67040;
  reg [31:0] p40_add_67680;
  reg [31:0] p40_add_67075;
  reg [31:0] p40_add_67850;
  reg [31:0] p40_add_67851;
  reg [31:0] p40_add_67213;
  reg [31:0] p40_add_67854;
  reg [31:0] p40_add_67536;
  reg [31:0] p40_add_67248;
  reg [31:0] p40_add_67705;
  reg [31:0] p40_add_67382;
  reg [31:0] p40_and_67855;
  reg [31:0] p40_add_67876;
  reg [31:0] p40_add_67417;
  reg [31:0] p40_add_67554;
  reg [31:0] p40_add_67589;
  reg [1:0] p40_bit_slice_67706;
  reg [31:0] p40_add_67724;
  reg [31:0] p40_add_67758;
  reg [31:0] p40_add_67894;
  reg [31:0] p40_add_67929;
  reg [31:0] p40_add_67946;
  always_ff @ (posedge clk) begin
    p40_add_65326 <= p39_add_65326;
    p40_add_66849 <= p39_add_66849;
    p40_add_66906 <= p39_add_66906;
    p40_add_67508 <= p39_add_67508;
    p40_add_67040 <= p39_add_67040;
    p40_add_67680 <= p39_add_67680;
    p40_add_67075 <= p39_add_67075;
    p40_add_67850 <= p40_add_67850_comb;
    p40_add_67851 <= p40_add_67851_comb;
    p40_add_67213 <= p39_add_67213;
    p40_add_67854 <= p40_add_67854_comb;
    p40_add_67536 <= p39_add_67536;
    p40_add_67248 <= p39_add_67248;
    p40_add_67705 <= p39_add_67705;
    p40_add_67382 <= p39_add_67382;
    p40_and_67855 <= p40_and_67855_comb;
    p40_add_67876 <= p40_add_67876_comb;
    p40_add_67417 <= p39_add_67417;
    p40_add_67554 <= p39_add_67554;
    p40_add_67589 <= p39_add_67589;
    p40_bit_slice_67706 <= p39_bit_slice_67706;
    p40_add_67724 <= p39_add_67724;
    p40_add_67758 <= p39_add_67758;
    p40_add_67894 <= p40_add_67894_comb;
    p40_add_67929 <= p40_add_67929_comb;
    p40_add_67946 <= p40_add_67946_comb;
  end

  // ===== Pipe stage 41:
  wire [31:0] p41_and_68026_comb;
  wire [31:0] p41_add_68020_comb;
  wire [31:0] p41_add_68021_comb;
  wire [31:0] p41_add_68024_comb;
  wire [31:0] p41_add_68045_comb;
  wire [31:0] p41_add_68064_comb;
  wire [31:0] p41_add_68098_comb;
  wire [31:0] p41_add_68099_comb;
  wire [31:0] p41_add_68022_comb;
  wire [31:0] p41_add_68025_comb;
  wire [31:0] p41_add_68047_comb;
  wire [31:0] p41_add_68065_comb;
  wire [31:0] p41_add_68100_comb;
  assign p41_and_68026_comb = p40_add_67876 & p40_add_67705;
  assign p41_add_68020_comb = {p40_add_67851[5:0] ^ p40_add_67851[10:5] ^ p40_add_67851[24:19], p40_add_67851[31:27] ^ p40_add_67851[4:0] ^ p40_add_67851[18:14], p40_add_67851[26:13] ^ p40_add_67851[31:18] ^ p40_add_67851[13:0], p40_add_67851[12:6] ^ p40_add_67851[17:11] ^ p40_add_67851[31:25]} + (p40_add_67851 & p40_add_67680 ^ ~(p40_add_67851 | ~p40_add_67508));
  assign p41_add_68021_comb = p41_add_68020_comb + p40_add_67854;
  assign p41_add_68024_comb = p40_add_67248 + 32'ha81a_664b;
  assign p41_add_68045_comb = (p41_and_68026_comb ^ p40_add_67876 & p40_add_67536 ^ p40_and_67855) + p40_add_67850;
  assign p41_add_68064_comb = p40_add_67417 + {p40_add_65326[6:4] ^ p40_add_65326[17:15], p40_add_65326[3:0] ^ p40_add_65326[14:11] ^ p40_add_65326[31:28], p40_add_65326[31:21] ^ p40_add_65326[10:0] ^ p40_add_65326[27:17], p40_add_65326[20:7] ^ p40_add_65326[31:18] ^ p40_add_65326[16:3]};
  assign p41_add_68098_comb = p40_add_67554 + {p40_add_66849[6:4] ^ p40_add_66849[17:15], p40_add_66849[3:0] ^ p40_add_66849[14:11] ^ p40_add_66849[31:28], p40_add_66849[31:21] ^ p40_add_66849[10:0] ^ p40_add_66849[27:17], p40_add_66849[20:7] ^ p40_add_66849[31:18] ^ p40_add_66849[16:3]};
  assign p41_add_68099_comb = {p40_add_67929[16:7] ^ p40_add_67929[18:9], p40_add_67929[6:0] ^ p40_add_67929[8:2] ^ p40_add_67929[31:25], p40_add_67929[31:30] ^ p40_add_67929[1:0] ^ p40_add_67929[24:23], p40_add_67929[29:17] ^ p40_add_67929[31:19] ^ p40_add_67929[22:10]} + p40_add_65326;
  assign p41_add_68022_comb = p41_add_68021_comb + p40_add_67536;
  assign p41_add_68025_comb = p40_add_67508 + p41_add_68024_comb;
  assign p41_add_68047_comb = p41_add_68045_comb + {p40_add_67876[1:0] ^ p40_add_67876[12:11] ^ p40_add_67876[21:20], p40_add_67876[31:21] ^ p40_add_67876[10:0] ^ p40_add_67876[19:9], p40_add_67876[20:12] ^ p40_add_67876[31:23] ^ p40_add_67876[8:0], p40_add_67876[11:2] ^ p40_add_67876[22:13] ^ p40_add_67876[31:22]};
  assign p41_add_68065_comb = p41_add_68064_comb + p40_add_67946;
  assign p41_add_68100_comb = p41_add_68098_comb + p41_add_68099_comb;

  // Registers for pipe stage 41:
  reg [31:0] p41_add_66849;
  reg [31:0] p41_add_66906;
  reg [31:0] p41_add_67040;
  reg [31:0] p41_add_67680;
  reg [31:0] p41_add_67075;
  reg [31:0] p41_add_67851;
  reg [31:0] p41_add_67213;
  reg [31:0] p41_add_68021;
  reg [31:0] p41_add_68022;
  reg [31:0] p41_add_67248;
  reg [31:0] p41_add_68025;
  reg [31:0] p41_add_67705;
  reg [31:0] p41_add_67382;
  reg [31:0] p41_add_67876;
  reg [31:0] p41_add_67417;
  reg [31:0] p41_and_68026;
  reg [31:0] p41_add_68047;
  reg [31:0] p41_add_67554;
  reg [31:0] p41_add_67589;
  reg [1:0] p41_bit_slice_67706;
  reg [31:0] p41_add_67724;
  reg [31:0] p41_add_67758;
  reg [31:0] p41_add_67894;
  reg [31:0] p41_add_67929;
  reg [31:0] p41_add_68065;
  reg [31:0] p41_add_68100;
  always_ff @ (posedge clk) begin
    p41_add_66849 <= p40_add_66849;
    p41_add_66906 <= p40_add_66906;
    p41_add_67040 <= p40_add_67040;
    p41_add_67680 <= p40_add_67680;
    p41_add_67075 <= p40_add_67075;
    p41_add_67851 <= p40_add_67851;
    p41_add_67213 <= p40_add_67213;
    p41_add_68021 <= p41_add_68021_comb;
    p41_add_68022 <= p41_add_68022_comb;
    p41_add_67248 <= p40_add_67248;
    p41_add_68025 <= p41_add_68025_comb;
    p41_add_67705 <= p40_add_67705;
    p41_add_67382 <= p40_add_67382;
    p41_add_67876 <= p40_add_67876;
    p41_add_67417 <= p40_add_67417;
    p41_and_68026 <= p41_and_68026_comb;
    p41_add_68047 <= p41_add_68047_comb;
    p41_add_67554 <= p40_add_67554;
    p41_add_67589 <= p40_add_67589;
    p41_bit_slice_67706 <= p40_bit_slice_67706;
    p41_add_67724 <= p40_add_67724;
    p41_add_67758 <= p40_add_67758;
    p41_add_67894 <= p40_add_67894;
    p41_add_67929 <= p40_add_67929;
    p41_add_68065 <= p41_add_68065_comb;
    p41_add_68100 <= p41_add_68100_comb;
  end

  // ===== Pipe stage 42:
  wire [1:0] p42_bit_slice_68205_comb;
  wire [31:0] p42_add_68237_comb;
  wire [31:0] p42_add_68238_comb;
  wire [31:0] p42_add_68239_comb;
  wire [31:0] p42_and_68183_comb;
  wire [31:0] p42_add_68174_comb;
  wire [27:0] p42_add_68179_comb;
  wire [31:0] p42_add_68175_comb;
  wire [31:0] p42_add_68202_comb;
  wire [31:0] p42_add_68272_comb;
  wire [31:0] p42_add_68273_comb;
  wire [31:0] p42_add_68176_comb;
  wire [31:0] p42_add_68182_comb;
  wire [31:0] p42_add_68204_comb;
  wire [31:0] p42_add_68274_comb;
  wire [31:0] p42_add_68291_comb;
  wire [3:0] p42_xor_68294_comb;
  assign p42_bit_slice_68205_comb = p41_add_68065[1:0];
  assign p42_add_68237_comb = p41_add_67589 + {p41_add_66906[6:4] ^ p41_add_66906[17:15], p41_add_66906[3:0] ^ p41_add_66906[14:11] ^ p41_add_66906[31:28], p41_add_66906[31:21] ^ p41_add_66906[10:0] ^ p41_add_66906[27:17], p41_add_66906[20:7] ^ p41_add_66906[31:18] ^ p41_add_66906[16:3]};
  assign p42_add_68238_comb = {p41_add_68065[16:7] ^ p41_add_68065[18:9], p41_add_68065[6:0] ^ p41_add_68065[8:2] ^ p41_add_68065[31:25], p41_add_68065[31:30] ^ p42_bit_slice_68205_comb ^ p41_add_68065[24:23], p41_add_68065[29:17] ^ p41_add_68065[31:19] ^ p41_add_68065[22:10]} + p41_add_66849;
  assign p42_add_68239_comb = p42_add_68237_comb + p42_add_68238_comb;
  assign p42_and_68183_comb = p41_add_68047 & p41_add_67876;
  assign p42_add_68174_comb = {p41_add_68022[5:0] ^ p41_add_68022[10:5] ^ p41_add_68022[24:19], p41_add_68022[31:27] ^ p41_add_68022[4:0] ^ p41_add_68022[18:14], p41_add_68022[26:13] ^ p41_add_68022[31:18] ^ p41_add_68022[13:0], p41_add_68022[12:6] ^ p41_add_68022[17:11] ^ p41_add_68022[31:25]} + (p41_add_68022 & p41_add_67851 ^ ~(p41_add_68022 | ~p41_add_67680));
  assign p42_add_68179_comb = p41_add_67382[31:4] + 28'hc24_b8b7;
  assign p42_add_68175_comb = p42_add_68174_comb + p41_add_68025;
  assign p42_add_68202_comb = (p42_and_68183_comb ^ p41_add_68047 & p41_add_67705 ^ p41_and_68026) + p41_add_68021;
  assign p42_add_68272_comb = p41_add_67724 + {p41_add_67040[6:4] ^ p41_add_67040[17:15], p41_add_67040[3:0] ^ p41_add_67040[14:11] ^ p41_add_67040[31:28], p41_add_67040[31:21] ^ p41_add_67040[10:0] ^ p41_add_67040[27:17], p41_add_67040[20:7] ^ p41_add_67040[31:18] ^ p41_add_67040[16:3]};
  assign p42_add_68273_comb = {p41_add_68100[16:7] ^ p41_add_68100[18:9], p41_add_68100[6:0] ^ p41_add_68100[8:2] ^ p41_add_68100[31:25], p41_add_68100[31:30] ^ p41_add_68100[1:0] ^ p41_add_68100[24:23], p41_add_68100[29:17] ^ p41_add_68100[31:19] ^ p41_add_68100[22:10]} + p41_add_66906;
  assign p42_add_68176_comb = p42_add_68175_comb + p41_add_67705;
  assign p42_add_68182_comb = {p42_add_68179_comb, p41_add_67382[3:0]} + p41_add_67680;
  assign p42_add_68204_comb = p42_add_68202_comb + {p41_add_68047[1:0] ^ p41_add_68047[12:11] ^ p41_add_68047[21:20], p41_add_68047[31:21] ^ p41_add_68047[10:0] ^ p41_add_68047[19:9], p41_add_68047[20:12] ^ p41_add_68047[31:23] ^ p41_add_68047[8:0], p41_add_68047[11:2] ^ p41_add_68047[22:13] ^ p41_add_68047[31:22]};
  assign p42_add_68274_comb = p42_add_68272_comb + p42_add_68273_comb;
  assign p42_add_68291_comb = {p42_add_68239_comb[16:7] ^ p42_add_68239_comb[18:9], p42_add_68239_comb[6:0] ^ p42_add_68239_comb[8:2] ^ p42_add_68239_comb[31:25], p42_add_68239_comb[31:30] ^ p42_add_68239_comb[1:0] ^ p42_add_68239_comb[24:23], p42_add_68239_comb[29:17] ^ p42_add_68239_comb[31:19] ^ p42_add_68239_comb[22:10]} + p41_add_67040;
  assign p42_xor_68294_comb = p41_add_67382[3:0] ^ p41_add_67382[14:11] ^ p41_add_67382[31:28];

  // Registers for pipe stage 42:
  reg [31:0] p42_add_67075;
  reg [31:0] p42_add_67851;
  reg [31:0] p42_add_67213;
  reg [31:0] p42_add_68022;
  reg [31:0] p42_add_67248;
  reg [31:0] p42_add_68175;
  reg [31:0] p42_add_68176;
  reg [31:0] p42_add_67382;
  reg [31:0] p42_add_68182;
  reg [31:0] p42_add_67876;
  reg [31:0] p42_add_67417;
  reg [31:0] p42_add_68047;
  reg [31:0] p42_add_67554;
  reg [31:0] p42_and_68183;
  reg [31:0] p42_add_68204;
  reg [31:0] p42_add_67589;
  reg [1:0] p42_bit_slice_67706;
  reg [31:0] p42_add_67724;
  reg [31:0] p42_add_67758;
  reg [31:0] p42_add_67894;
  reg [31:0] p42_add_67929;
  reg [31:0] p42_add_68065;
  reg [1:0] p42_bit_slice_68205;
  reg [31:0] p42_add_68100;
  reg [31:0] p42_add_68239;
  reg [31:0] p42_add_68274;
  reg [31:0] p42_add_68291;
  reg [3:0] p42_xor_68294;
  always_ff @ (posedge clk) begin
    p42_add_67075 <= p41_add_67075;
    p42_add_67851 <= p41_add_67851;
    p42_add_67213 <= p41_add_67213;
    p42_add_68022 <= p41_add_68022;
    p42_add_67248 <= p41_add_67248;
    p42_add_68175 <= p42_add_68175_comb;
    p42_add_68176 <= p42_add_68176_comb;
    p42_add_67382 <= p41_add_67382;
    p42_add_68182 <= p42_add_68182_comb;
    p42_add_67876 <= p41_add_67876;
    p42_add_67417 <= p41_add_67417;
    p42_add_68047 <= p41_add_68047;
    p42_add_67554 <= p41_add_67554;
    p42_and_68183 <= p42_and_68183_comb;
    p42_add_68204 <= p42_add_68204_comb;
    p42_add_67589 <= p41_add_67589;
    p42_bit_slice_67706 <= p41_bit_slice_67706;
    p42_add_67724 <= p41_add_67724;
    p42_add_67758 <= p41_add_67758;
    p42_add_67894 <= p41_add_67894;
    p42_add_67929 <= p41_add_67929;
    p42_add_68065 <= p41_add_68065;
    p42_bit_slice_68205 <= p42_bit_slice_68205_comb;
    p42_add_68100 <= p41_add_68100;
    p42_add_68239 <= p42_add_68239_comb;
    p42_add_68274 <= p42_add_68274_comb;
    p42_add_68291 <= p42_add_68291_comb;
    p42_xor_68294 <= p42_xor_68294_comb;
  end

  // ===== Pipe stage 43:
  wire [31:0] p43_add_68416_comb;
  wire [31:0] p43_add_68417_comb;
  wire [31:0] p43_and_68378_comb;
  wire [31:0] p43_add_68372_comb;
  wire [31:0] p43_add_68373_comb;
  wire [31:0] p43_add_68376_comb;
  wire [31:0] p43_add_68397_comb;
  wire [31:0] p43_add_68450_comb;
  wire [31:0] p43_add_68451_comb;
  wire [31:0] p43_add_68374_comb;
  wire [31:0] p43_add_68377_comb;
  wire [31:0] p43_add_68399_comb;
  wire [31:0] p43_add_68452_comb;
  wire [31:0] p43_add_68469_comb;
  assign p43_add_68416_comb = p42_add_67758 + {p42_add_67075[6:4] ^ p42_add_67075[17:15], p42_add_67075[3:0] ^ p42_add_67075[14:11] ^ p42_add_67075[31:28], p42_add_67075[31:21] ^ p42_add_67075[10:0] ^ p42_add_67075[27:17], p42_add_67075[20:7] ^ p42_add_67075[31:18] ^ p42_add_67075[16:3]};
  assign p43_add_68417_comb = p43_add_68416_comb + p42_add_68291;
  assign p43_and_68378_comb = p42_add_68204 & p42_add_68047;
  assign p43_add_68372_comb = (p42_add_68176 & p42_add_68022 ^ ~(p42_add_68176 | ~p42_add_67851)) + {p42_add_68176[5:0] ^ p42_add_68176[10:5] ^ p42_add_68176[24:19], p42_add_68176[31:27] ^ p42_add_68176[4:0] ^ p42_add_68176[18:14], p42_add_68176[26:13] ^ p42_add_68176[31:18] ^ p42_add_68176[13:0], p42_add_68176[12:6] ^ p42_add_68176[17:11] ^ p42_add_68176[31:25]};
  assign p43_add_68373_comb = p43_add_68372_comb + p42_add_68182;
  assign p43_add_68376_comb = p42_add_67417 + 32'hc76c_51a3;
  assign p43_add_68397_comb = (p43_and_68378_comb ^ p42_add_68204 & p42_add_67876 ^ p42_and_68183) + p42_add_68175;
  assign p43_add_68450_comb = p42_add_67894 + {p42_add_67213[6:4] ^ p42_add_67213[17:15], p42_add_67213[3:0] ^ p42_add_67213[14:11] ^ p42_add_67213[31:28], p42_add_67213[31:21] ^ p42_add_67213[10:0] ^ p42_add_67213[27:17], p42_add_67213[20:7] ^ p42_add_67213[31:18] ^ p42_add_67213[16:3]};
  assign p43_add_68451_comb = {p42_add_68274[16:7] ^ p42_add_68274[18:9], p42_add_68274[6:0] ^ p42_add_68274[8:2] ^ p42_add_68274[31:25], p42_add_68274[31:30] ^ p42_add_68274[1:0] ^ p42_add_68274[24:23], p42_add_68274[29:17] ^ p42_add_68274[31:19] ^ p42_add_68274[22:10]} + p42_add_67075;
  assign p43_add_68374_comb = p43_add_68373_comb + p42_add_67876;
  assign p43_add_68377_comb = p42_add_67851 + p43_add_68376_comb;
  assign p43_add_68399_comb = p43_add_68397_comb + {p42_add_68204[1:0] ^ p42_add_68204[12:11] ^ p42_add_68204[21:20], p42_add_68204[31:21] ^ p42_add_68204[10:0] ^ p42_add_68204[19:9], p42_add_68204[20:12] ^ p42_add_68204[31:23] ^ p42_add_68204[8:0], p42_add_68204[11:2] ^ p42_add_68204[22:13] ^ p42_add_68204[31:22]};
  assign p43_add_68452_comb = p43_add_68450_comb + p43_add_68451_comb;
  assign p43_add_68469_comb = {p43_add_68417_comb[16:7] ^ p43_add_68417_comb[18:9], p43_add_68417_comb[6:0] ^ p43_add_68417_comb[8:2] ^ p43_add_68417_comb[31:25], p43_add_68417_comb[31:30] ^ p43_add_68417_comb[1:0] ^ p43_add_68417_comb[24:23], p43_add_68417_comb[29:17] ^ p43_add_68417_comb[31:19] ^ p43_add_68417_comb[22:10]} + p42_add_67213;

  // Registers for pipe stage 43:
  reg [31:0] p43_add_68022;
  reg [31:0] p43_add_67248;
  reg [31:0] p43_add_68176;
  reg [31:0] p43_add_67382;
  reg [31:0] p43_add_68373;
  reg [31:0] p43_add_68374;
  reg [31:0] p43_add_67417;
  reg [31:0] p43_add_68377;
  reg [31:0] p43_add_68047;
  reg [31:0] p43_add_67554;
  reg [31:0] p43_add_68204;
  reg [31:0] p43_add_67589;
  reg [1:0] p43_bit_slice_67706;
  reg [31:0] p43_and_68378;
  reg [31:0] p43_add_68399;
  reg [31:0] p43_add_67724;
  reg [31:0] p43_add_67758;
  reg [31:0] p43_add_67894;
  reg [31:0] p43_add_67929;
  reg [31:0] p43_add_68065;
  reg [1:0] p43_bit_slice_68205;
  reg [31:0] p43_add_68100;
  reg [31:0] p43_add_68239;
  reg [31:0] p43_add_68274;
  reg [31:0] p43_add_68417;
  reg [31:0] p43_add_68452;
  reg [31:0] p43_add_68469;
  reg [3:0] p43_xor_68294;
  always_ff @ (posedge clk) begin
    p43_add_68022 <= p42_add_68022;
    p43_add_67248 <= p42_add_67248;
    p43_add_68176 <= p42_add_68176;
    p43_add_67382 <= p42_add_67382;
    p43_add_68373 <= p43_add_68373_comb;
    p43_add_68374 <= p43_add_68374_comb;
    p43_add_67417 <= p42_add_67417;
    p43_add_68377 <= p43_add_68377_comb;
    p43_add_68047 <= p42_add_68047;
    p43_add_67554 <= p42_add_67554;
    p43_add_68204 <= p42_add_68204;
    p43_add_67589 <= p42_add_67589;
    p43_bit_slice_67706 <= p42_bit_slice_67706;
    p43_and_68378 <= p43_and_68378_comb;
    p43_add_68399 <= p43_add_68399_comb;
    p43_add_67724 <= p42_add_67724;
    p43_add_67758 <= p42_add_67758;
    p43_add_67894 <= p42_add_67894;
    p43_add_67929 <= p42_add_67929;
    p43_add_68065 <= p42_add_68065;
    p43_bit_slice_68205 <= p42_bit_slice_68205;
    p43_add_68100 <= p42_add_68100;
    p43_add_68239 <= p42_add_68239;
    p43_add_68274 <= p42_add_68274;
    p43_add_68417 <= p43_add_68417_comb;
    p43_add_68452 <= p43_add_68452_comb;
    p43_add_68469 <= p43_add_68469_comb;
    p43_xor_68294 <= p42_xor_68294;
  end

  // ===== Pipe stage 44:
  wire [31:0] p44_add_68600_comb;
  wire [31:0] p44_add_68601_comb;
  wire [31:0] p44_and_68553_comb;
  wire [31:0] p44_add_68547_comb;
  wire [31:0] p44_add_68548_comb;
  wire [31:0] p44_add_68551_comb;
  wire [31:0] p44_add_68572_comb;
  wire [28:0] p44_add_68577_comb;
  wire [29:0] p44_add_68582_comb;
  wire [31:0] p44_add_68630_comb;
  wire [31:0] p44_add_68631_comb;
  wire [31:0] p44_add_68549_comb;
  wire [31:0] p44_add_68552_comb;
  wire [31:0] p44_add_68574_comb;
  wire [31:0] p44_concat_68579_comb;
  wire [31:0] p44_concat_68583_comb;
  wire [31:0] p44_add_68632_comb;
  wire [31:0] p44_add_68649_comb;
  assign p44_add_68600_comb = p43_add_67929 + {p43_add_67248[6:4] ^ p43_add_67248[17:15], p43_add_67248[3:0] ^ p43_add_67248[14:11] ^ p43_add_67248[31:28], p43_add_67248[31:21] ^ p43_add_67248[10:0] ^ p43_add_67248[27:17], p43_add_67248[20:7] ^ p43_add_67248[31:18] ^ p43_add_67248[16:3]};
  assign p44_add_68601_comb = p44_add_68600_comb + p43_add_68469;
  assign p44_and_68553_comb = p43_add_68399 & p43_add_68204;
  assign p44_add_68547_comb = {p43_add_68374[5:0] ^ p43_add_68374[10:5] ^ p43_add_68374[24:19], p43_add_68374[31:27] ^ p43_add_68374[4:0] ^ p43_add_68374[18:14], p43_add_68374[26:13] ^ p43_add_68374[31:18] ^ p43_add_68374[13:0], p43_add_68374[12:6] ^ p43_add_68374[17:11] ^ p43_add_68374[31:25]} + (p43_add_68374 & p43_add_68176 ^ ~(p43_add_68374 | ~p43_add_68022));
  assign p44_add_68548_comb = p44_add_68547_comb + p43_add_68377;
  assign p44_add_68551_comb = p43_add_67554 + 32'hd192_e819;
  assign p44_add_68572_comb = (p44_and_68553_comb ^ p43_add_68399 & p43_add_68047 ^ p43_and_68378) + p43_add_68373;
  assign p44_add_68577_comb = p43_add_67929[31:3] + 29'h03c6_ed81;
  assign p44_add_68582_comb = p43_add_68065[31:2] + 30'h09d2_1dd3;
  assign p44_add_68630_comb = p43_add_68065 + {p43_add_67382[6:4] ^ p43_add_67382[17:15], p43_xor_68294, p43_add_67382[31:21] ^ p43_add_67382[10:0] ^ p43_add_67382[27:17], p43_add_67382[20:7] ^ p43_add_67382[31:18] ^ p43_add_67382[16:3]};
  assign p44_add_68631_comb = {p43_add_68452[16:7] ^ p43_add_68452[18:9], p43_add_68452[6:0] ^ p43_add_68452[8:2] ^ p43_add_68452[31:25], p43_add_68452[31:30] ^ p43_add_68452[1:0] ^ p43_add_68452[24:23], p43_add_68452[29:17] ^ p43_add_68452[31:19] ^ p43_add_68452[22:10]} + p43_add_67248;
  assign p44_add_68549_comb = p44_add_68548_comb + p43_add_68047;
  assign p44_add_68552_comb = p43_add_68022 + p44_add_68551_comb;
  assign p44_add_68574_comb = p44_add_68572_comb + {p43_add_68399[1:0] ^ p43_add_68399[12:11] ^ p43_add_68399[21:20], p43_add_68399[31:21] ^ p43_add_68399[10:0] ^ p43_add_68399[19:9], p43_add_68399[20:12] ^ p43_add_68399[31:23] ^ p43_add_68399[8:0], p43_add_68399[11:2] ^ p43_add_68399[22:13] ^ p43_add_68399[31:22]};
  assign p44_concat_68579_comb = {p44_add_68577_comb, p43_add_67929[2:0]};
  assign p44_concat_68583_comb = {p44_add_68582_comb, p43_bit_slice_68205};
  assign p44_add_68632_comb = p44_add_68630_comb + p44_add_68631_comb;
  assign p44_add_68649_comb = {p44_add_68601_comb[16:7] ^ p44_add_68601_comb[18:9], p44_add_68601_comb[6:0] ^ p44_add_68601_comb[8:2] ^ p44_add_68601_comb[31:25], p44_add_68601_comb[31:30] ^ p44_add_68601_comb[1:0] ^ p44_add_68601_comb[24:23], p44_add_68601_comb[29:17] ^ p44_add_68601_comb[31:19] ^ p44_add_68601_comb[22:10]} + p43_add_67382;

  // Registers for pipe stage 44:
  reg [31:0] p44_add_68176;
  reg [31:0] p44_add_68374;
  reg [31:0] p44_add_67417;
  reg [31:0] p44_add_68548;
  reg [31:0] p44_add_68549;
  reg [31:0] p44_add_67554;
  reg [31:0] p44_add_68552;
  reg [31:0] p44_add_68204;
  reg [31:0] p44_add_67589;
  reg [1:0] p44_bit_slice_67706;
  reg [31:0] p44_add_68399;
  reg [31:0] p44_add_67724;
  reg [31:0] p44_and_68553;
  reg [31:0] p44_add_68574;
  reg [31:0] p44_add_67758;
  reg [31:0] p44_add_67894;
  reg [31:0] p44_concat_68579;
  reg [31:0] p44_concat_68583;
  reg [31:0] p44_add_68100;
  reg [31:0] p44_add_68239;
  reg [31:0] p44_add_68274;
  reg [31:0] p44_add_68417;
  reg [31:0] p44_add_68452;
  reg [31:0] p44_add_68601;
  reg [31:0] p44_add_68632;
  reg [31:0] p44_add_68649;
  always_ff @ (posedge clk) begin
    p44_add_68176 <= p43_add_68176;
    p44_add_68374 <= p43_add_68374;
    p44_add_67417 <= p43_add_67417;
    p44_add_68548 <= p44_add_68548_comb;
    p44_add_68549 <= p44_add_68549_comb;
    p44_add_67554 <= p43_add_67554;
    p44_add_68552 <= p44_add_68552_comb;
    p44_add_68204 <= p43_add_68204;
    p44_add_67589 <= p43_add_67589;
    p44_bit_slice_67706 <= p43_bit_slice_67706;
    p44_add_68399 <= p43_add_68399;
    p44_add_67724 <= p43_add_67724;
    p44_and_68553 <= p44_and_68553_comb;
    p44_add_68574 <= p44_add_68574_comb;
    p44_add_67758 <= p43_add_67758;
    p44_add_67894 <= p43_add_67894;
    p44_concat_68579 <= p44_concat_68579_comb;
    p44_concat_68583 <= p44_concat_68583_comb;
    p44_add_68100 <= p43_add_68100;
    p44_add_68239 <= p43_add_68239;
    p44_add_68274 <= p43_add_68274;
    p44_add_68417 <= p43_add_68417;
    p44_add_68452 <= p43_add_68452;
    p44_add_68601 <= p44_add_68601_comb;
    p44_add_68632 <= p44_add_68632_comb;
    p44_add_68649 <= p44_add_68649_comb;
  end

  // ===== Pipe stage 45:
  wire [31:0] p45_add_68775_comb;
  wire [31:0] p45_add_68776_comb;
  wire [31:0] p45_and_68731_comb;
  wire [31:0] p45_add_68723_comb;
  wire [29:0] p45_add_68728_comb;
  wire [31:0] p45_add_68724_comb;
  wire [31:0] p45_add_68750_comb;
  wire [29:0] p45_add_68779_comb;
  wire [31:0] p45_add_68814_comb;
  wire [31:0] p45_add_68815_comb;
  wire [31:0] p45_add_68725_comb;
  wire [31:0] p45_add_68730_comb;
  wire [31:0] p45_add_68752_comb;
  wire [31:0] p45_add_68754_comb;
  wire [31:0] p45_add_68756_comb;
  wire [31:0] p45_add_68769_comb;
  wire [31:0] p45_concat_68803_comb;
  wire [31:0] p45_add_68816_comb;
  wire [31:0] p45_add_68832_comb;
  assign p45_add_68775_comb = p44_add_68100 + {p44_add_67417[6:4] ^ p44_add_67417[17:15], p44_add_67417[3:0] ^ p44_add_67417[14:11] ^ p44_add_67417[31:28], p44_add_67417[31:21] ^ p44_add_67417[10:0] ^ p44_add_67417[27:17], p44_add_67417[20:7] ^ p44_add_67417[31:18] ^ p44_add_67417[16:3]};
  assign p45_add_68776_comb = p45_add_68775_comb + p44_add_68649;
  assign p45_and_68731_comb = p44_add_68574 & p44_add_68399;
  assign p45_add_68723_comb = {p44_add_68549[5:0] ^ p44_add_68549[10:5] ^ p44_add_68549[24:19], p44_add_68549[31:27] ^ p44_add_68549[4:0] ^ p44_add_68549[18:14], p44_add_68549[26:13] ^ p44_add_68549[31:18] ^ p44_add_68549[13:0], p44_add_68549[12:6] ^ p44_add_68549[17:11] ^ p44_add_68549[31:25]} + (p44_add_68549 & p44_add_68374 ^ ~(p44_add_68549 | ~p44_add_68176));
  assign p45_add_68728_comb = p44_add_67589[31:2] + 30'h35a6_4189;
  assign p45_add_68724_comb = p45_add_68723_comb + p44_add_68552;
  assign p45_add_68750_comb = (p45_and_68731_comb ^ p44_add_68574 & p44_add_68204 ^ p44_and_68553) + p44_add_68548;
  assign p45_add_68779_comb = p45_add_68776_comb[31:2] + 30'h2132_1e05;
  assign p45_add_68814_comb = p44_add_68239 + {p44_add_67554[6:4] ^ p44_add_67554[17:15], p44_add_67554[3:0] ^ p44_add_67554[14:11] ^ p44_add_67554[31:28], p44_add_67554[31:21] ^ p44_add_67554[10:0] ^ p44_add_67554[27:17], p44_add_67554[20:7] ^ p44_add_67554[31:18] ^ p44_add_67554[16:3]};
  assign p45_add_68815_comb = {p44_add_68632[16:7] ^ p44_add_68632[18:9], p44_add_68632[6:0] ^ p44_add_68632[8:2] ^ p44_add_68632[31:25], p44_add_68632[31:30] ^ p44_add_68632[1:0] ^ p44_add_68632[24:23], p44_add_68632[29:17] ^ p44_add_68632[31:19] ^ p44_add_68632[22:10]} + p44_add_67417;
  assign p45_add_68725_comb = p45_add_68724_comb + p44_add_68204;
  assign p45_add_68730_comb = {p45_add_68728_comb, p44_bit_slice_67706} + p44_add_68176;
  assign p45_add_68752_comb = p45_add_68750_comb + {p44_add_68574[1:0] ^ p44_add_68574[12:11] ^ p44_add_68574[21:20], p44_add_68574[31:21] ^ p44_add_68574[10:0] ^ p44_add_68574[19:9], p44_add_68574[20:12] ^ p44_add_68574[31:23] ^ p44_add_68574[8:0], p44_add_68574[11:2] ^ p44_add_68574[22:13] ^ p44_add_68574[31:22]};
  assign p45_add_68754_comb = p44_add_68100 + 32'h34b0_bcb5;
  assign p45_add_68756_comb = p44_add_68239 + 32'h391c_0cb3;
  assign p45_add_68769_comb = p44_add_68632 + 32'h78a5_636f;
  assign p45_concat_68803_comb = {p45_add_68779_comb, p45_add_68776_comb[1:0]};
  assign p45_add_68816_comb = p45_add_68814_comb + p45_add_68815_comb;
  assign p45_add_68832_comb = {p45_add_68776_comb[16:7] ^ p45_add_68776_comb[18:9], p45_add_68776_comb[6:0] ^ p45_add_68776_comb[8:2] ^ p45_add_68776_comb[31:25], p45_add_68776_comb[31:30] ^ p45_add_68776_comb[1:0] ^ p45_add_68776_comb[24:23], p45_add_68776_comb[29:17] ^ p45_add_68776_comb[31:19] ^ p45_add_68776_comb[22:10]} + p44_add_67554;

  // Registers for pipe stage 45:
  reg [31:0] p45_add_68374;
  reg [31:0] p45_add_68549;
  reg [31:0] p45_add_68724;
  reg [31:0] p45_add_68725;
  reg [31:0] p45_add_67589;
  reg [31:0] p45_add_68730;
  reg [31:0] p45_add_68399;
  reg [31:0] p45_add_67724;
  reg [31:0] p45_add_68574;
  reg [31:0] p45_add_67758;
  reg [31:0] p45_and_68731;
  reg [31:0] p45_add_68752;
  reg [31:0] p45_add_67894;
  reg [31:0] p45_concat_68579;
  reg [31:0] p45_concat_68583;
  reg [31:0] p45_add_68754;
  reg [31:0] p45_add_68756;
  reg [31:0] p45_add_68274;
  reg [31:0] p45_add_68417;
  reg [31:0] p45_add_68452;
  reg [31:0] p45_add_68601;
  reg [31:0] p45_add_68769;
  reg [31:0] p45_concat_68803;
  reg [31:0] p45_add_68816;
  reg [31:0] p45_add_68832;
  always_ff @ (posedge clk) begin
    p45_add_68374 <= p44_add_68374;
    p45_add_68549 <= p44_add_68549;
    p45_add_68724 <= p45_add_68724_comb;
    p45_add_68725 <= p45_add_68725_comb;
    p45_add_67589 <= p44_add_67589;
    p45_add_68730 <= p45_add_68730_comb;
    p45_add_68399 <= p44_add_68399;
    p45_add_67724 <= p44_add_67724;
    p45_add_68574 <= p44_add_68574;
    p45_add_67758 <= p44_add_67758;
    p45_and_68731 <= p45_and_68731_comb;
    p45_add_68752 <= p45_add_68752_comb;
    p45_add_67894 <= p44_add_67894;
    p45_concat_68579 <= p44_concat_68579;
    p45_concat_68583 <= p44_concat_68583;
    p45_add_68754 <= p45_add_68754_comb;
    p45_add_68756 <= p45_add_68756_comb;
    p45_add_68274 <= p44_add_68274;
    p45_add_68417 <= p44_add_68417;
    p45_add_68452 <= p44_add_68452;
    p45_add_68601 <= p44_add_68601;
    p45_add_68769 <= p45_add_68769_comb;
    p45_concat_68803 <= p45_concat_68803_comb;
    p45_add_68816 <= p45_add_68816_comb;
    p45_add_68832 <= p45_add_68832_comb;
  end

  // ===== Pipe stage 46:
  wire [31:0] p46_and_68910_comb;
  wire [31:0] p46_add_68904_comb;
  wire [31:0] p46_add_68905_comb;
  wire [31:0] p46_add_68908_comb;
  wire [31:0] p46_add_68929_comb;
  wire [30:0] p46_add_68934_comb;
  wire [28:0] p46_add_68941_comb;
  wire [31:0] p46_add_68960_comb;
  wire [31:0] p46_add_68994_comb;
  wire [31:0] p46_add_68995_comb;
  wire [31:0] p46_add_68906_comb;
  wire [31:0] p46_add_68909_comb;
  wire [31:0] p46_add_68931_comb;
  wire [31:0] p46_concat_68936_comb;
  wire [31:0] p46_add_68938_comb;
  wire [31:0] p46_concat_68954_comb;
  wire [31:0] p46_add_68961_comb;
  wire [31:0] p46_add_68996_comb;
  assign p46_and_68910_comb = p45_add_68752 & p45_add_68574;
  assign p46_add_68904_comb = (p45_add_68725 & p45_add_68549 ^ ~(p45_add_68725 | ~p45_add_68374)) + {p45_add_68725[5:0] ^ p45_add_68725[10:5] ^ p45_add_68725[24:19], p45_add_68725[31:27] ^ p45_add_68725[4:0] ^ p45_add_68725[18:14], p45_add_68725[26:13] ^ p45_add_68725[31:18] ^ p45_add_68725[13:0], p45_add_68725[12:6] ^ p45_add_68725[17:11] ^ p45_add_68725[31:25]};
  assign p46_add_68905_comb = p46_add_68904_comb + p45_add_68730;
  assign p46_add_68908_comb = p45_add_67724 + 32'hf40e_3585;
  assign p46_add_68929_comb = (p46_and_68910_comb ^ p45_add_68752 & p45_add_68399 ^ p45_and_68731) + p45_add_68724;
  assign p46_add_68934_comb = p45_add_68274[31:1] + 31'h276c_5525;
  assign p46_add_68941_comb = p45_add_68816[31:3] + 29'h1198_e041;
  assign p46_add_68960_comb = p45_add_68274 + {p45_add_67589[6:4] ^ p45_add_67589[17:15], p45_add_67589[3:0] ^ p45_add_67589[14:11] ^ p45_add_67589[31:28], p45_add_67589[31:21] ^ p45_add_67589[10:0] ^ p45_add_67589[27:17], p45_add_67589[20:7] ^ p45_add_67589[31:18] ^ p45_add_67589[16:3]};
  assign p46_add_68994_comb = p45_add_68417 + {p45_add_67724[6:4] ^ p45_add_67724[17:15], p45_add_67724[3:0] ^ p45_add_67724[14:11] ^ p45_add_67724[31:28], p45_add_67724[31:21] ^ p45_add_67724[10:0] ^ p45_add_67724[27:17], p45_add_67724[20:7] ^ p45_add_67724[31:18] ^ p45_add_67724[16:3]};
  assign p46_add_68995_comb = {p45_add_68816[16:7] ^ p45_add_68816[18:9], p45_add_68816[6:0] ^ p45_add_68816[8:2] ^ p45_add_68816[31:25], p45_add_68816[31:30] ^ p45_add_68816[1:0] ^ p45_add_68816[24:23], p45_add_68816[29:17] ^ p45_add_68816[31:19] ^ p45_add_68816[22:10]} + p45_add_67589;
  assign p46_add_68906_comb = p46_add_68905_comb + p45_add_68399;
  assign p46_add_68909_comb = p45_add_68374 + p46_add_68908_comb;
  assign p46_add_68931_comb = p46_add_68929_comb + {p45_add_68752[1:0] ^ p45_add_68752[12:11] ^ p45_add_68752[21:20], p45_add_68752[31:21] ^ p45_add_68752[10:0] ^ p45_add_68752[19:9], p45_add_68752[20:12] ^ p45_add_68752[31:23] ^ p45_add_68752[8:0], p45_add_68752[11:2] ^ p45_add_68752[22:13] ^ p45_add_68752[31:22]};
  assign p46_concat_68936_comb = {p46_add_68934_comb, p45_add_68274[0]};
  assign p46_add_68938_comb = p45_add_68417 + 32'h5b9c_ca4f;
  assign p46_concat_68954_comb = {p46_add_68941_comb, p45_add_68816[2:0]};
  assign p46_add_68961_comb = p46_add_68960_comb + p45_add_68832;
  assign p46_add_68996_comb = p46_add_68994_comb + p46_add_68995_comb;

  // Registers for pipe stage 46:
  reg [31:0] p46_add_68549;
  reg [31:0] p46_add_68725;
  reg [31:0] p46_add_68905;
  reg [31:0] p46_add_68906;
  reg [31:0] p46_add_67724;
  reg [31:0] p46_add_68909;
  reg [31:0] p46_add_68574;
  reg [31:0] p46_add_67758;
  reg [31:0] p46_add_68752;
  reg [31:0] p46_add_67894;
  reg [31:0] p46_and_68910;
  reg [31:0] p46_add_68931;
  reg [31:0] p46_concat_68579;
  reg [31:0] p46_concat_68583;
  reg [31:0] p46_add_68754;
  reg [31:0] p46_add_68756;
  reg [31:0] p46_concat_68936;
  reg [31:0] p46_add_68938;
  reg [31:0] p46_add_68452;
  reg [31:0] p46_add_68601;
  reg [31:0] p46_add_68769;
  reg [31:0] p46_concat_68803;
  reg [31:0] p46_concat_68954;
  reg [31:0] p46_add_68961;
  reg [31:0] p46_add_68996;
  always_ff @ (posedge clk) begin
    p46_add_68549 <= p45_add_68549;
    p46_add_68725 <= p45_add_68725;
    p46_add_68905 <= p46_add_68905_comb;
    p46_add_68906 <= p46_add_68906_comb;
    p46_add_67724 <= p45_add_67724;
    p46_add_68909 <= p46_add_68909_comb;
    p46_add_68574 <= p45_add_68574;
    p46_add_67758 <= p45_add_67758;
    p46_add_68752 <= p45_add_68752;
    p46_add_67894 <= p45_add_67894;
    p46_and_68910 <= p46_and_68910_comb;
    p46_add_68931 <= p46_add_68931_comb;
    p46_concat_68579 <= p45_concat_68579;
    p46_concat_68583 <= p45_concat_68583;
    p46_add_68754 <= p45_add_68754;
    p46_add_68756 <= p45_add_68756;
    p46_concat_68936 <= p46_concat_68936_comb;
    p46_add_68938 <= p46_add_68938_comb;
    p46_add_68452 <= p45_add_68452;
    p46_add_68601 <= p45_add_68601;
    p46_add_68769 <= p45_add_68769;
    p46_concat_68803 <= p45_concat_68803;
    p46_concat_68954 <= p46_concat_68954_comb;
    p46_add_68961 <= p46_add_68961_comb;
    p46_add_68996 <= p46_add_68996_comb;
  end

  // ===== Pipe stage 47:
  wire [31:0] p47_and_69077_comb;
  wire [31:0] p47_add_69068_comb;
  wire [27:0] p47_add_69073_comb;
  wire [31:0] p47_add_69069_comb;
  wire [31:0] p47_add_69097_comb;
  wire [31:0] p47_add_69070_comb;
  wire [31:0] p47_add_69076_comb;
  wire [31:0] p47_add_69096_comb;
  wire [31:0] p47_add_69099_comb;
  wire [3:0] p47_xor_69102_comb;
  assign p47_and_69077_comb = p46_add_68931 & p46_add_68752;
  assign p47_add_69068_comb = {p46_add_68906[5:0] ^ p46_add_68906[10:5] ^ p46_add_68906[24:19], p46_add_68906[31:27] ^ p46_add_68906[4:0] ^ p46_add_68906[18:14], p46_add_68906[26:13] ^ p46_add_68906[31:18] ^ p46_add_68906[13:0], p46_add_68906[12:6] ^ p46_add_68906[17:11] ^ p46_add_68906[31:25]} + (p46_add_68906 & p46_add_68725 ^ ~(p46_add_68906 | ~p46_add_68549));
  assign p47_add_69073_comb = p46_add_67758[31:4] + 28'h106_aa07;
  assign p47_add_69069_comb = p47_add_69068_comb + p46_add_68909;
  assign p47_add_69097_comb = (p47_and_69077_comb ^ p46_add_68931 & p46_add_68574 ^ p46_and_68910) + p46_add_68905;
  assign p47_add_69070_comb = p47_add_69069_comb + p46_add_68574;
  assign p47_add_69076_comb = {p47_add_69073_comb, p46_add_67758[3:0]} + p46_add_68549;
  assign p47_add_69096_comb = p46_concat_68579 + p46_add_68906;
  assign p47_add_69099_comb = p47_add_69097_comb + {p46_add_68931[1:0] ^ p46_add_68931[12:11] ^ p46_add_68931[21:20], p46_add_68931[31:21] ^ p46_add_68931[10:0] ^ p46_add_68931[19:9], p46_add_68931[20:12] ^ p46_add_68931[31:23] ^ p46_add_68931[8:0], p46_add_68931[11:2] ^ p46_add_68931[22:13] ^ p46_add_68931[31:22]};
  assign p47_xor_69102_comb = p46_add_67758[3:0] ^ p46_add_67758[14:11] ^ p46_add_67758[31:28];

  // Registers for pipe stage 47:
  reg [31:0] p47_add_68725;
  reg [31:0] p47_add_68906;
  reg [31:0] p47_add_67724;
  reg [31:0] p47_add_69069;
  reg [31:0] p47_add_69070;
  reg [31:0] p47_add_67758;
  reg [31:0] p47_add_69076;
  reg [31:0] p47_add_68752;
  reg [31:0] p47_add_67894;
  reg [31:0] p47_add_68931;
  reg [31:0] p47_and_69077;
  reg [31:0] p47_add_69096;
  reg [31:0] p47_add_69099;
  reg [31:0] p47_concat_68583;
  reg [31:0] p47_add_68754;
  reg [31:0] p47_add_68756;
  reg [31:0] p47_concat_68936;
  reg [31:0] p47_add_68938;
  reg [31:0] p47_add_68452;
  reg [31:0] p47_add_68601;
  reg [31:0] p47_add_68769;
  reg [31:0] p47_concat_68803;
  reg [31:0] p47_concat_68954;
  reg [31:0] p47_add_68961;
  reg [31:0] p47_add_68996;
  reg [3:0] p47_xor_69102;
  always_ff @ (posedge clk) begin
    p47_add_68725 <= p46_add_68725;
    p47_add_68906 <= p46_add_68906;
    p47_add_67724 <= p46_add_67724;
    p47_add_69069 <= p47_add_69069_comb;
    p47_add_69070 <= p47_add_69070_comb;
    p47_add_67758 <= p46_add_67758;
    p47_add_69076 <= p47_add_69076_comb;
    p47_add_68752 <= p46_add_68752;
    p47_add_67894 <= p46_add_67894;
    p47_add_68931 <= p46_add_68931;
    p47_and_69077 <= p47_and_69077_comb;
    p47_add_69096 <= p47_add_69096_comb;
    p47_add_69099 <= p47_add_69099_comb;
    p47_concat_68583 <= p46_concat_68583;
    p47_add_68754 <= p46_add_68754;
    p47_add_68756 <= p46_add_68756;
    p47_concat_68936 <= p46_concat_68936;
    p47_add_68938 <= p46_add_68938;
    p47_add_68452 <= p46_add_68452;
    p47_add_68601 <= p46_add_68601;
    p47_add_68769 <= p46_add_68769;
    p47_concat_68803 <= p46_concat_68803;
    p47_concat_68954 <= p46_concat_68954;
    p47_add_68961 <= p46_add_68961;
    p47_add_68996 <= p46_add_68996;
    p47_xor_69102 <= p47_xor_69102_comb;
  end

  // ===== Pipe stage 48:
  wire [12:0] p48_xor_69228_comb;
  wire [31:0] p48_add_69176_comb;
  wire [31:0] p48_and_69187_comb;
  wire [31:0] p48_add_69177_comb;
  wire [30:0] p48_add_69183_comb;
  wire [30:0] p48_add_69251_comb;
  wire [31:0] p48_add_69178_comb;
  wire [31:0] p48_add_69207_comb;
  wire [30:0] p48_add_69212_comb;
  wire [31:0] p48_add_69253_comb;
  wire [31:0] p48_nor_69182_comb;
  wire [31:0] p48_add_69186_comb;
  wire [31:0] p48_add_69206_comb;
  wire [31:0] p48_add_69209_comb;
  wire [31:0] p48_concat_69214_comb;
  wire [31:0] p48_add_69216_comb;
  wire [31:0] p48_add_69255_comb;
  assign p48_xor_69228_comb = p47_add_68996[29:17] ^ p47_add_68996[31:19] ^ p47_add_68996[22:10];
  assign p48_add_69176_comb = (p47_add_69070 & p47_add_68906 ^ ~(p47_add_69070 | ~p47_add_68725)) + {p47_add_69070[5:0] ^ p47_add_69070[10:5] ^ p47_add_69070[24:19], p47_add_69070[31:27] ^ p47_add_69070[4:0] ^ p47_add_69070[18:14], p47_add_69070[26:13] ^ p47_add_69070[31:18] ^ p47_add_69070[13:0], p47_add_69070[12:6] ^ p47_add_69070[17:11] ^ p47_add_69070[31:25]};
  assign p48_and_69187_comb = p47_add_69099 & p47_add_68931;
  assign p48_add_69177_comb = p48_add_69176_comb + p47_add_69076;
  assign p48_add_69183_comb = p47_add_67894[31:1] + 31'h0cd2_608b;
  assign p48_add_69251_comb = {p47_add_68996[16:7] ^ p47_add_68996[18:9], p47_add_68996[6:0] ^ p47_add_68996[8:2] ^ p47_add_68996[31:25], p47_add_68996[31:30] ^ p47_add_68996[1:0] ^ p47_add_68996[24:23], p48_xor_69228_comb[12:1]} + 31'h6338_bc79;
  assign p48_add_69178_comb = p48_add_69177_comb + p47_add_68752;
  assign p48_add_69207_comb = (p48_and_69187_comb ^ p47_add_69099 & p47_add_68752 ^ p47_and_69077) + p47_add_69069;
  assign p48_add_69212_comb = p47_add_68601[31:1] + 31'h3a47_c177;
  assign p48_add_69253_comb = {p47_add_67894[6:4] ^ p47_add_67894[17:15], p47_add_67894[3:0] ^ p47_add_67894[14:11] ^ p47_add_67894[31:28], p47_add_67894[31:21] ^ p47_add_67894[10:0] ^ p47_add_67894[27:17], p47_add_67894[20:7] ^ p47_add_67894[31:18] ^ p47_add_67894[16:3]} + p47_add_68601;
  assign p48_nor_69182_comb = ~(p48_add_69178_comb | ~p47_add_68906);
  assign p48_add_69186_comb = {p48_add_69183_comb, p47_add_67894[0]} + p47_add_68725;
  assign p48_add_69206_comb = p47_concat_68583 + p47_add_69070;
  assign p48_add_69209_comb = p48_add_69207_comb + {p47_add_69099[1:0] ^ p47_add_69099[12:11] ^ p47_add_69099[21:20], p47_add_69099[31:21] ^ p47_add_69099[10:0] ^ p47_add_69099[19:9], p47_add_69099[20:12] ^ p47_add_69099[31:23] ^ p47_add_69099[8:0], p47_add_69099[11:2] ^ p47_add_69099[22:13] ^ p47_add_69099[31:22]};
  assign p48_concat_69214_comb = {p48_add_69212_comb, p47_add_68601[0]};
  assign p48_add_69216_comb = p47_add_68996 + 32'ha450_6ceb;
  assign p48_add_69255_comb = p48_add_69253_comb + {p48_add_69251_comb, p48_xor_69228_comb[0]};

  // Registers for pipe stage 48:
  reg [31:0] p48_add_67724;
  reg [31:0] p48_add_69070;
  reg [31:0] p48_add_67758;
  reg [31:0] p48_add_69177;
  reg [31:0] p48_add_69178;
  reg [31:0] p48_nor_69182;
  reg [31:0] p48_add_69186;
  reg [31:0] p48_add_68931;
  reg [31:0] p48_add_69096;
  reg [31:0] p48_add_69099;
  reg [31:0] p48_and_69187;
  reg [31:0] p48_add_69206;
  reg [31:0] p48_add_69209;
  reg [31:0] p48_add_68754;
  reg [31:0] p48_add_68756;
  reg [31:0] p48_concat_68936;
  reg [31:0] p48_add_68938;
  reg [31:0] p48_add_68452;
  reg [31:0] p48_concat_69214;
  reg [31:0] p48_add_68769;
  reg [31:0] p48_concat_68803;
  reg [31:0] p48_concat_68954;
  reg [31:0] p48_add_68961;
  reg [31:0] p48_add_69216;
  reg [3:0] p48_xor_69102;
  reg [31:0] p48_add_69255;
  always_ff @ (posedge clk) begin
    p48_add_67724 <= p47_add_67724;
    p48_add_69070 <= p47_add_69070;
    p48_add_67758 <= p47_add_67758;
    p48_add_69177 <= p48_add_69177_comb;
    p48_add_69178 <= p48_add_69178_comb;
    p48_nor_69182 <= p48_nor_69182_comb;
    p48_add_69186 <= p48_add_69186_comb;
    p48_add_68931 <= p47_add_68931;
    p48_add_69096 <= p47_add_69096;
    p48_add_69099 <= p47_add_69099;
    p48_and_69187 <= p48_and_69187_comb;
    p48_add_69206 <= p48_add_69206_comb;
    p48_add_69209 <= p48_add_69209_comb;
    p48_add_68754 <= p47_add_68754;
    p48_add_68756 <= p47_add_68756;
    p48_concat_68936 <= p47_concat_68936;
    p48_add_68938 <= p47_add_68938;
    p48_add_68452 <= p47_add_68452;
    p48_concat_69214 <= p48_concat_69214_comb;
    p48_add_68769 <= p47_add_68769;
    p48_concat_68803 <= p47_concat_68803;
    p48_concat_68954 <= p47_concat_68954;
    p48_add_68961 <= p47_add_68961;
    p48_add_69216 <= p48_add_69216_comb;
    p48_xor_69102 <= p47_xor_69102;
    p48_add_69255 <= p48_add_69255_comb;
  end

  // ===== Pipe stage 49:
  wire [31:0] p49_add_69327_comb;
  wire [31:0] p49_and_69332_comb;
  wire [31:0] p49_add_69328_comb;
  wire [31:0] p49_add_69329_comb;
  wire [31:0] p49_add_69352_comb;
  wire [31:0] p49_nor_69331_comb;
  wire [31:0] p49_add_69351_comb;
  wire [31:0] p49_add_69354_comb;
  assign p49_add_69327_comb = (p48_add_69178 & p48_add_69070 ^ p48_nor_69182) + {p48_add_69178[5:0] ^ p48_add_69178[10:5] ^ p48_add_69178[24:19], p48_add_69178[31:27] ^ p48_add_69178[4:0] ^ p48_add_69178[18:14], p48_add_69178[26:13] ^ p48_add_69178[31:18] ^ p48_add_69178[13:0], p48_add_69178[12:6] ^ p48_add_69178[17:11] ^ p48_add_69178[31:25]};
  assign p49_and_69332_comb = p48_add_69209 & p48_add_69099;
  assign p49_add_69328_comb = p49_add_69327_comb + p48_add_69186;
  assign p49_add_69329_comb = p49_add_69328_comb + p48_add_68931;
  assign p49_add_69352_comb = (p49_and_69332_comb ^ p48_add_69209 & p48_add_68931 ^ p48_and_69187) + p48_add_69177;
  assign p49_nor_69331_comb = ~(p49_add_69329_comb | ~p48_add_69070);
  assign p49_add_69351_comb = p48_add_69178 + p48_add_68754;
  assign p49_add_69354_comb = p49_add_69352_comb + {p48_add_69209[1:0] ^ p48_add_69209[12:11] ^ p48_add_69209[21:20], p48_add_69209[31:21] ^ p48_add_69209[10:0] ^ p48_add_69209[19:9], p48_add_69209[20:12] ^ p48_add_69209[31:23] ^ p48_add_69209[8:0], p48_add_69209[11:2] ^ p48_add_69209[22:13] ^ p48_add_69209[31:22]};

  // Registers for pipe stage 49:
  reg [31:0] p49_add_67724;
  reg [31:0] p49_add_67758;
  reg [31:0] p49_add_69178;
  reg [31:0] p49_add_69328;
  reg [31:0] p49_add_69329;
  reg [31:0] p49_nor_69331;
  reg [31:0] p49_add_69096;
  reg [31:0] p49_add_69099;
  reg [31:0] p49_add_69206;
  reg [31:0] p49_add_69209;
  reg [31:0] p49_and_69332;
  reg [31:0] p49_add_69351;
  reg [31:0] p49_add_69354;
  reg [31:0] p49_add_68756;
  reg [31:0] p49_concat_68936;
  reg [31:0] p49_add_68938;
  reg [31:0] p49_add_68452;
  reg [31:0] p49_concat_69214;
  reg [31:0] p49_add_68769;
  reg [31:0] p49_concat_68803;
  reg [31:0] p49_concat_68954;
  reg [31:0] p49_add_68961;
  reg [31:0] p49_add_69216;
  reg [3:0] p49_xor_69102;
  reg [31:0] p49_add_69255;
  always_ff @ (posedge clk) begin
    p49_add_67724 <= p48_add_67724;
    p49_add_67758 <= p48_add_67758;
    p49_add_69178 <= p48_add_69178;
    p49_add_69328 <= p49_add_69328_comb;
    p49_add_69329 <= p49_add_69329_comb;
    p49_nor_69331 <= p49_nor_69331_comb;
    p49_add_69096 <= p48_add_69096;
    p49_add_69099 <= p48_add_69099;
    p49_add_69206 <= p48_add_69206;
    p49_add_69209 <= p48_add_69209;
    p49_and_69332 <= p49_and_69332_comb;
    p49_add_69351 <= p49_add_69351_comb;
    p49_add_69354 <= p49_add_69354_comb;
    p49_add_68756 <= p48_add_68756;
    p49_concat_68936 <= p48_concat_68936;
    p49_add_68938 <= p48_add_68938;
    p49_add_68452 <= p48_add_68452;
    p49_concat_69214 <= p48_concat_69214;
    p49_add_68769 <= p48_add_68769;
    p49_concat_68803 <= p48_concat_68803;
    p49_concat_68954 <= p48_concat_68954;
    p49_add_68961 <= p48_add_68961;
    p49_add_69216 <= p48_add_69216;
    p49_xor_69102 <= p48_xor_69102;
    p49_add_69255 <= p48_add_69255;
  end

  // ===== Pipe stage 50:
  wire [31:0] p50_add_69424_comb;
  wire [31:0] p50_and_69429_comb;
  wire [31:0] p50_add_69425_comb;
  wire [31:0] p50_add_69426_comb;
  wire [31:0] p50_add_69449_comb;
  wire [31:0] p50_nor_69428_comb;
  wire [31:0] p50_add_69448_comb;
  wire [31:0] p50_add_69451_comb;
  assign p50_add_69424_comb = (p49_add_69329 & p49_add_69178 ^ p49_nor_69331) + {p49_add_69329[5:0] ^ p49_add_69329[10:5] ^ p49_add_69329[24:19], p49_add_69329[31:27] ^ p49_add_69329[4:0] ^ p49_add_69329[18:14], p49_add_69329[26:13] ^ p49_add_69329[31:18] ^ p49_add_69329[13:0], p49_add_69329[12:6] ^ p49_add_69329[17:11] ^ p49_add_69329[31:25]};
  assign p50_and_69429_comb = p49_add_69354 & p49_add_69209;
  assign p50_add_69425_comb = p50_add_69424_comb + p49_add_69096;
  assign p50_add_69426_comb = p50_add_69425_comb + p49_add_69099;
  assign p50_add_69449_comb = (p50_and_69429_comb ^ p49_add_69354 & p49_add_69099 ^ p49_and_69332) + p49_add_69328;
  assign p50_nor_69428_comb = ~(p50_add_69426_comb | ~p49_add_69178);
  assign p50_add_69448_comb = p49_add_69329 + p49_add_68756;
  assign p50_add_69451_comb = p50_add_69449_comb + {p49_add_69354[1:0] ^ p49_add_69354[12:11] ^ p49_add_69354[21:20], p49_add_69354[31:21] ^ p49_add_69354[10:0] ^ p49_add_69354[19:9], p49_add_69354[20:12] ^ p49_add_69354[31:23] ^ p49_add_69354[8:0], p49_add_69354[11:2] ^ p49_add_69354[22:13] ^ p49_add_69354[31:22]};

  // Registers for pipe stage 50:
  reg [31:0] p50_add_67724;
  reg [31:0] p50_add_67758;
  reg [31:0] p50_add_69329;
  reg [31:0] p50_add_69425;
  reg [31:0] p50_add_69426;
  reg [31:0] p50_nor_69428;
  reg [31:0] p50_add_69206;
  reg [31:0] p50_add_69209;
  reg [31:0] p50_add_69351;
  reg [31:0] p50_add_69354;
  reg [31:0] p50_and_69429;
  reg [31:0] p50_add_69448;
  reg [31:0] p50_add_69451;
  reg [31:0] p50_concat_68936;
  reg [31:0] p50_add_68938;
  reg [31:0] p50_add_68452;
  reg [31:0] p50_concat_69214;
  reg [31:0] p50_add_68769;
  reg [31:0] p50_concat_68803;
  reg [31:0] p50_concat_68954;
  reg [31:0] p50_add_68961;
  reg [31:0] p50_add_69216;
  reg [3:0] p50_xor_69102;
  reg [31:0] p50_add_69255;
  always_ff @ (posedge clk) begin
    p50_add_67724 <= p49_add_67724;
    p50_add_67758 <= p49_add_67758;
    p50_add_69329 <= p49_add_69329;
    p50_add_69425 <= p50_add_69425_comb;
    p50_add_69426 <= p50_add_69426_comb;
    p50_nor_69428 <= p50_nor_69428_comb;
    p50_add_69206 <= p49_add_69206;
    p50_add_69209 <= p49_add_69209;
    p50_add_69351 <= p49_add_69351;
    p50_add_69354 <= p49_add_69354;
    p50_and_69429 <= p50_and_69429_comb;
    p50_add_69448 <= p50_add_69448_comb;
    p50_add_69451 <= p50_add_69451_comb;
    p50_concat_68936 <= p49_concat_68936;
    p50_add_68938 <= p49_add_68938;
    p50_add_68452 <= p49_add_68452;
    p50_concat_69214 <= p49_concat_69214;
    p50_add_68769 <= p49_add_68769;
    p50_concat_68803 <= p49_concat_68803;
    p50_concat_68954 <= p49_concat_68954;
    p50_add_68961 <= p49_add_68961;
    p50_add_69216 <= p49_add_69216;
    p50_xor_69102 <= p49_xor_69102;
    p50_add_69255 <= p49_add_69255;
  end

  // ===== Pipe stage 51:
  wire [31:0] p51_add_69519_comb;
  wire [31:0] p51_and_69524_comb;
  wire [31:0] p51_add_69520_comb;
  wire [31:0] p51_add_69521_comb;
  wire [31:0] p51_add_69544_comb;
  wire [31:0] p51_nor_69523_comb;
  wire [31:0] p51_add_69543_comb;
  wire [31:0] p51_add_69546_comb;
  assign p51_add_69519_comb = (p50_add_69426 & p50_add_69329 ^ p50_nor_69428) + {p50_add_69426[5:0] ^ p50_add_69426[10:5] ^ p50_add_69426[24:19], p50_add_69426[31:27] ^ p50_add_69426[4:0] ^ p50_add_69426[18:14], p50_add_69426[26:13] ^ p50_add_69426[31:18] ^ p50_add_69426[13:0], p50_add_69426[12:6] ^ p50_add_69426[17:11] ^ p50_add_69426[31:25]};
  assign p51_and_69524_comb = p50_add_69451 & p50_add_69354;
  assign p51_add_69520_comb = p51_add_69519_comb + p50_add_69206;
  assign p51_add_69521_comb = p51_add_69520_comb + p50_add_69209;
  assign p51_add_69544_comb = (p51_and_69524_comb ^ p50_add_69451 & p50_add_69209 ^ p50_and_69429) + p50_add_69425;
  assign p51_nor_69523_comb = ~(p51_add_69521_comb | ~p50_add_69329);
  assign p51_add_69543_comb = p50_concat_68936 + p50_add_69426;
  assign p51_add_69546_comb = p51_add_69544_comb + {p50_add_69451[1:0] ^ p50_add_69451[12:11] ^ p50_add_69451[21:20], p50_add_69451[31:21] ^ p50_add_69451[10:0] ^ p50_add_69451[19:9], p50_add_69451[20:12] ^ p50_add_69451[31:23] ^ p50_add_69451[8:0], p50_add_69451[11:2] ^ p50_add_69451[22:13] ^ p50_add_69451[31:22]};

  // Registers for pipe stage 51:
  reg [31:0] p51_add_67724;
  reg [31:0] p51_add_67758;
  reg [31:0] p51_add_69426;
  reg [31:0] p51_add_69520;
  reg [31:0] p51_add_69521;
  reg [31:0] p51_nor_69523;
  reg [31:0] p51_add_69351;
  reg [31:0] p51_add_69354;
  reg [31:0] p51_add_69448;
  reg [31:0] p51_add_69451;
  reg [31:0] p51_and_69524;
  reg [31:0] p51_add_69543;
  reg [31:0] p51_add_69546;
  reg [31:0] p51_add_68938;
  reg [31:0] p51_add_68452;
  reg [31:0] p51_concat_69214;
  reg [31:0] p51_add_68769;
  reg [31:0] p51_concat_68803;
  reg [31:0] p51_concat_68954;
  reg [31:0] p51_add_68961;
  reg [31:0] p51_add_69216;
  reg [3:0] p51_xor_69102;
  reg [31:0] p51_add_69255;
  always_ff @ (posedge clk) begin
    p51_add_67724 <= p50_add_67724;
    p51_add_67758 <= p50_add_67758;
    p51_add_69426 <= p50_add_69426;
    p51_add_69520 <= p51_add_69520_comb;
    p51_add_69521 <= p51_add_69521_comb;
    p51_nor_69523 <= p51_nor_69523_comb;
    p51_add_69351 <= p50_add_69351;
    p51_add_69354 <= p50_add_69354;
    p51_add_69448 <= p50_add_69448;
    p51_add_69451 <= p50_add_69451;
    p51_and_69524 <= p51_and_69524_comb;
    p51_add_69543 <= p51_add_69543_comb;
    p51_add_69546 <= p51_add_69546_comb;
    p51_add_68938 <= p50_add_68938;
    p51_add_68452 <= p50_add_68452;
    p51_concat_69214 <= p50_concat_69214;
    p51_add_68769 <= p50_add_68769;
    p51_concat_68803 <= p50_concat_68803;
    p51_concat_68954 <= p50_concat_68954;
    p51_add_68961 <= p50_add_68961;
    p51_add_69216 <= p50_add_69216;
    p51_xor_69102 <= p50_xor_69102;
    p51_add_69255 <= p50_add_69255;
  end

  // ===== Pipe stage 52:
  wire [31:0] p52_add_69612_comb;
  wire [31:0] p52_and_69617_comb;
  wire [31:0] p52_add_69613_comb;
  wire [31:0] p52_add_69614_comb;
  wire [31:0] p52_add_69637_comb;
  wire [31:0] p52_nor_69616_comb;
  wire [31:0] p52_add_69636_comb;
  wire [31:0] p52_add_69639_comb;
  assign p52_add_69612_comb = {p51_add_69521[5:0] ^ p51_add_69521[10:5] ^ p51_add_69521[24:19], p51_add_69521[31:27] ^ p51_add_69521[4:0] ^ p51_add_69521[18:14], p51_add_69521[26:13] ^ p51_add_69521[31:18] ^ p51_add_69521[13:0], p51_add_69521[12:6] ^ p51_add_69521[17:11] ^ p51_add_69521[31:25]} + (p51_add_69521 & p51_add_69426 ^ p51_nor_69523);
  assign p52_and_69617_comb = p51_add_69546 & p51_add_69451;
  assign p52_add_69613_comb = p52_add_69612_comb + p51_add_69351;
  assign p52_add_69614_comb = p52_add_69613_comb + p51_add_69354;
  assign p52_add_69637_comb = (p52_and_69617_comb ^ p51_add_69546 & p51_add_69354 ^ p51_and_69524) + p51_add_69520;
  assign p52_nor_69616_comb = ~(p52_add_69614_comb | ~p51_add_69426);
  assign p52_add_69636_comb = p51_add_69521 + p51_add_68938;
  assign p52_add_69639_comb = p52_add_69637_comb + {p51_add_69546[1:0] ^ p51_add_69546[12:11] ^ p51_add_69546[21:20], p51_add_69546[31:21] ^ p51_add_69546[10:0] ^ p51_add_69546[19:9], p51_add_69546[20:12] ^ p51_add_69546[31:23] ^ p51_add_69546[8:0], p51_add_69546[11:2] ^ p51_add_69546[22:13] ^ p51_add_69546[31:22]};

  // Registers for pipe stage 52:
  reg [31:0] p52_add_67724;
  reg [31:0] p52_add_67758;
  reg [31:0] p52_add_69521;
  reg [31:0] p52_add_69613;
  reg [31:0] p52_add_69614;
  reg [31:0] p52_nor_69616;
  reg [31:0] p52_add_69448;
  reg [31:0] p52_add_69451;
  reg [31:0] p52_add_69543;
  reg [31:0] p52_add_69546;
  reg [31:0] p52_and_69617;
  reg [31:0] p52_add_69636;
  reg [31:0] p52_add_69639;
  reg [31:0] p52_add_68452;
  reg [31:0] p52_concat_69214;
  reg [31:0] p52_add_68769;
  reg [31:0] p52_concat_68803;
  reg [31:0] p52_concat_68954;
  reg [31:0] p52_add_68961;
  reg [31:0] p52_add_69216;
  reg [3:0] p52_xor_69102;
  reg [31:0] p52_add_69255;
  always_ff @ (posedge clk) begin
    p52_add_67724 <= p51_add_67724;
    p52_add_67758 <= p51_add_67758;
    p52_add_69521 <= p51_add_69521;
    p52_add_69613 <= p52_add_69613_comb;
    p52_add_69614 <= p52_add_69614_comb;
    p52_nor_69616 <= p52_nor_69616_comb;
    p52_add_69448 <= p51_add_69448;
    p52_add_69451 <= p51_add_69451;
    p52_add_69543 <= p51_add_69543;
    p52_add_69546 <= p51_add_69546;
    p52_and_69617 <= p52_and_69617_comb;
    p52_add_69636 <= p52_add_69636_comb;
    p52_add_69639 <= p52_add_69639_comb;
    p52_add_68452 <= p51_add_68452;
    p52_concat_69214 <= p51_concat_69214;
    p52_add_68769 <= p51_add_68769;
    p52_concat_68803 <= p51_concat_68803;
    p52_concat_68954 <= p51_concat_68954;
    p52_add_68961 <= p51_add_68961;
    p52_add_69216 <= p51_add_69216;
    p52_xor_69102 <= p51_xor_69102;
    p52_add_69255 <= p51_add_69255;
  end

  // ===== Pipe stage 53:
  wire [31:0] p53_add_69703_comb;
  wire [31:0] p53_and_69708_comb;
  wire [31:0] p53_add_69704_comb;
  wire [31:0] p53_add_69705_comb;
  wire [31:0] p53_add_69727_comb;
  wire [31:0] p53_nor_69707_comb;
  wire [31:0] p53_add_69729_comb;
  assign p53_add_69703_comb = {p52_add_69614[5:0] ^ p52_add_69614[10:5] ^ p52_add_69614[24:19], p52_add_69614[31:27] ^ p52_add_69614[4:0] ^ p52_add_69614[18:14], p52_add_69614[26:13] ^ p52_add_69614[31:18] ^ p52_add_69614[13:0], p52_add_69614[12:6] ^ p52_add_69614[17:11] ^ p52_add_69614[31:25]} + (p52_add_69614 & p52_add_69521 ^ p52_nor_69616);
  assign p53_and_69708_comb = p52_add_69639 & p52_add_69546;
  assign p53_add_69704_comb = p53_add_69703_comb + p52_add_69448;
  assign p53_add_69705_comb = p53_add_69704_comb + p52_add_69451;
  assign p53_add_69727_comb = (p53_and_69708_comb ^ p52_add_69639 & p52_add_69451 ^ p52_and_69617) + p52_add_69613;
  assign p53_nor_69707_comb = ~(p53_add_69705_comb | ~p52_add_69521);
  assign p53_add_69729_comb = p53_add_69727_comb + {p52_add_69639[1:0] ^ p52_add_69639[12:11] ^ p52_add_69639[21:20], p52_add_69639[31:21] ^ p52_add_69639[10:0] ^ p52_add_69639[19:9], p52_add_69639[20:12] ^ p52_add_69639[31:23] ^ p52_add_69639[8:0], p52_add_69639[11:2] ^ p52_add_69639[22:13] ^ p52_add_69639[31:22]};

  // Registers for pipe stage 53:
  reg [31:0] p53_add_67724;
  reg [31:0] p53_add_67758;
  reg [31:0] p53_add_69614;
  reg [31:0] p53_add_69704;
  reg [31:0] p53_add_69705;
  reg [31:0] p53_nor_69707;
  reg [31:0] p53_add_69543;
  reg [31:0] p53_add_69546;
  reg [31:0] p53_add_69636;
  reg [31:0] p53_add_69639;
  reg [31:0] p53_add_68452;
  reg [31:0] p53_and_69708;
  reg [31:0] p53_add_69729;
  reg [31:0] p53_concat_69214;
  reg [31:0] p53_add_68769;
  reg [31:0] p53_concat_68803;
  reg [31:0] p53_concat_68954;
  reg [31:0] p53_add_68961;
  reg [31:0] p53_add_69216;
  reg [3:0] p53_xor_69102;
  reg [31:0] p53_add_69255;
  always_ff @ (posedge clk) begin
    p53_add_67724 <= p52_add_67724;
    p53_add_67758 <= p52_add_67758;
    p53_add_69614 <= p52_add_69614;
    p53_add_69704 <= p53_add_69704_comb;
    p53_add_69705 <= p53_add_69705_comb;
    p53_nor_69707 <= p53_nor_69707_comb;
    p53_add_69543 <= p52_add_69543;
    p53_add_69546 <= p52_add_69546;
    p53_add_69636 <= p52_add_69636;
    p53_add_69639 <= p52_add_69639;
    p53_add_68452 <= p52_add_68452;
    p53_and_69708 <= p53_and_69708_comb;
    p53_add_69729 <= p53_add_69729_comb;
    p53_concat_69214 <= p52_concat_69214;
    p53_add_68769 <= p52_add_68769;
    p53_concat_68803 <= p52_concat_68803;
    p53_concat_68954 <= p52_concat_68954;
    p53_add_68961 <= p52_add_68961;
    p53_add_69216 <= p52_add_69216;
    p53_xor_69102 <= p52_xor_69102;
    p53_add_69255 <= p52_add_69255;
  end

  // ===== Pipe stage 54:
  wire [31:0] p54_and_69794_comb;
  wire [31:0] p54_add_69791_comb;
  wire [31:0] p54_add_69792_comb;
  wire [31:0] p54_add_69814_comb;
  wire [31:0] p54_add_69793_comb;
  wire [31:0] p54_add_69813_comb;
  wire [31:0] p54_add_69816_comb;
  assign p54_and_69794_comb = p53_add_69729 & p53_add_69639;
  assign p54_add_69791_comb = (p53_add_69705 & p53_add_69614 ^ p53_nor_69707) + {p53_add_69705[5:0] ^ p53_add_69705[10:5] ^ p53_add_69705[24:19], p53_add_69705[31:27] ^ p53_add_69705[4:0] ^ p53_add_69705[18:14], p53_add_69705[26:13] ^ p53_add_69705[31:18] ^ p53_add_69705[13:0], p53_add_69705[12:6] ^ p53_add_69705[17:11] ^ p53_add_69705[31:25]};
  assign p54_add_69792_comb = p54_add_69791_comb + p53_add_69543;
  assign p54_add_69814_comb = (p54_and_69794_comb ^ p53_add_69729 & p53_add_69546 ^ p53_and_69708) + p53_add_69704;
  assign p54_add_69793_comb = p54_add_69792_comb + p53_add_69546;
  assign p54_add_69813_comb = p53_concat_69214 + p53_add_69705;
  assign p54_add_69816_comb = p54_add_69814_comb + {p53_add_69729[1:0] ^ p53_add_69729[12:11] ^ p53_add_69729[21:20], p53_add_69729[31:21] ^ p53_add_69729[10:0] ^ p53_add_69729[19:9], p53_add_69729[20:12] ^ p53_add_69729[31:23] ^ p53_add_69729[8:0], p53_add_69729[11:2] ^ p53_add_69729[22:13] ^ p53_add_69729[31:22]};

  // Registers for pipe stage 54:
  reg [31:0] p54_add_67724;
  reg [31:0] p54_add_67758;
  reg [31:0] p54_add_69614;
  reg [31:0] p54_add_69705;
  reg [31:0] p54_add_69792;
  reg [31:0] p54_add_69793;
  reg [31:0] p54_add_69636;
  reg [31:0] p54_add_69639;
  reg [31:0] p54_add_68452;
  reg [31:0] p54_add_69729;
  reg [31:0] p54_and_69794;
  reg [31:0] p54_add_69813;
  reg [31:0] p54_add_69816;
  reg [31:0] p54_add_68769;
  reg [31:0] p54_concat_68803;
  reg [31:0] p54_concat_68954;
  reg [31:0] p54_add_68961;
  reg [31:0] p54_add_69216;
  reg [3:0] p54_xor_69102;
  reg [31:0] p54_add_69255;
  always_ff @ (posedge clk) begin
    p54_add_67724 <= p53_add_67724;
    p54_add_67758 <= p53_add_67758;
    p54_add_69614 <= p53_add_69614;
    p54_add_69705 <= p53_add_69705;
    p54_add_69792 <= p54_add_69792_comb;
    p54_add_69793 <= p54_add_69793_comb;
    p54_add_69636 <= p53_add_69636;
    p54_add_69639 <= p53_add_69639;
    p54_add_68452 <= p53_add_68452;
    p54_add_69729 <= p53_add_69729;
    p54_and_69794 <= p54_and_69794_comb;
    p54_add_69813 <= p54_add_69813_comb;
    p54_add_69816 <= p54_add_69816_comb;
    p54_add_68769 <= p53_add_68769;
    p54_concat_68803 <= p53_concat_68803;
    p54_concat_68954 <= p53_concat_68954;
    p54_add_68961 <= p53_add_68961;
    p54_add_69216 <= p53_add_69216;
    p54_xor_69102 <= p53_xor_69102;
    p54_add_69255 <= p53_add_69255;
  end

  // ===== Pipe stage 55:
  wire [31:0] p55_add_69878_comb;
  wire [31:0] p55_and_69886_comb;
  wire [31:0] p55_add_69879_comb;
  wire [31:0] p55_add_69880_comb;
  wire [31:0] p55_add_69884_comb;
  wire [31:0] p55_add_69905_comb;
  wire [30:0] p55_add_69911_comb;
  wire [31:0] p55_add_69943_comb;
  wire [31:0] p55_add_69944_comb;
  wire [31:0] p55_nor_69882_comb;
  wire [31:0] p55_add_69885_comb;
  wire [31:0] p55_add_69907_comb;
  wire [31:0] p55_add_69908_comb;
  wire [31:0] p55_concat_69913_comb;
  wire [31:0] p55_add_69945_comb;
  assign p55_add_69878_comb = {p54_add_69793[5:0] ^ p54_add_69793[10:5] ^ p54_add_69793[24:19], p54_add_69793[31:27] ^ p54_add_69793[4:0] ^ p54_add_69793[18:14], p54_add_69793[26:13] ^ p54_add_69793[31:18] ^ p54_add_69793[13:0], p54_add_69793[12:6] ^ p54_add_69793[17:11] ^ p54_add_69793[31:25]} + (p54_add_69793 & p54_add_69705 ^ ~(p54_add_69793 | ~p54_add_69614));
  assign p55_and_69886_comb = p54_add_69816 & p54_add_69729;
  assign p55_add_69879_comb = p55_add_69878_comb + p54_add_69636;
  assign p55_add_69880_comb = p55_add_69879_comb + p54_add_69639;
  assign p55_add_69884_comb = p54_add_68452 + 32'h682e_6ff3;
  assign p55_add_69905_comb = (p55_and_69886_comb ^ p54_add_69816 & p54_add_69639 ^ p54_and_69794) + p54_add_69792;
  assign p55_add_69911_comb = p54_add_68961[31:1] + 31'h485f_7ffd;
  assign p55_add_69943_comb = {p54_add_67758[6:4] ^ p54_add_67758[17:15], p54_xor_69102, p54_add_67758[31:21] ^ p54_add_67758[10:0] ^ p54_add_67758[27:17], p54_add_67758[20:7] ^ p54_add_67758[31:18] ^ p54_add_67758[16:3]} + p54_add_68452;
  assign p55_add_69944_comb = {p54_add_68961[16:7] ^ p54_add_68961[18:9], p54_add_68961[6:0] ^ p54_add_68961[8:2] ^ p54_add_68961[31:25], p54_add_68961[31:30] ^ p54_add_68961[1:0] ^ p54_add_68961[24:23], p54_add_68961[29:17] ^ p54_add_68961[31:19] ^ p54_add_68961[22:10]} + 32'hbef9_a3f7;
  assign p55_nor_69882_comb = ~(p55_add_69880_comb | ~p54_add_69705);
  assign p55_add_69885_comb = p54_add_69614 + p55_add_69884_comb;
  assign p55_add_69907_comb = p55_add_69905_comb + {p54_add_69816[1:0] ^ p54_add_69816[12:11] ^ p54_add_69816[21:20], p54_add_69816[31:21] ^ p54_add_69816[10:0] ^ p54_add_69816[19:9], p54_add_69816[20:12] ^ p54_add_69816[31:23] ^ p54_add_69816[8:0], p54_add_69816[11:2] ^ p54_add_69816[22:13] ^ p54_add_69816[31:22]};
  assign p55_add_69908_comb = p54_add_69793 + p54_add_68769;
  assign p55_concat_69913_comb = {p55_add_69911_comb, p54_add_68961[0]};
  assign p55_add_69945_comb = p55_add_69943_comb + p55_add_69944_comb;

  // Registers for pipe stage 55:
  reg [31:0] p55_add_67724;
  reg [31:0] p55_add_67758;
  reg [31:0] p55_add_69793;
  reg [31:0] p55_add_69879;
  reg [31:0] p55_add_69880;
  reg [31:0] p55_nor_69882;
  reg [31:0] p55_add_69885;
  reg [31:0] p55_add_69729;
  reg [31:0] p55_add_69813;
  reg [31:0] p55_add_69816;
  reg [31:0] p55_and_69886;
  reg [31:0] p55_add_69907;
  reg [31:0] p55_add_69908;
  reg [31:0] p55_concat_68803;
  reg [31:0] p55_concat_68954;
  reg [31:0] p55_concat_69913;
  reg [31:0] p55_add_69216;
  reg [31:0] p55_add_69255;
  reg [31:0] p55_add_69945;
  always_ff @ (posedge clk) begin
    p55_add_67724 <= p54_add_67724;
    p55_add_67758 <= p54_add_67758;
    p55_add_69793 <= p54_add_69793;
    p55_add_69879 <= p55_add_69879_comb;
    p55_add_69880 <= p55_add_69880_comb;
    p55_nor_69882 <= p55_nor_69882_comb;
    p55_add_69885 <= p55_add_69885_comb;
    p55_add_69729 <= p54_add_69729;
    p55_add_69813 <= p54_add_69813;
    p55_add_69816 <= p54_add_69816;
    p55_and_69886 <= p55_and_69886_comb;
    p55_add_69907 <= p55_add_69907_comb;
    p55_add_69908 <= p55_add_69908_comb;
    p55_concat_68803 <= p54_concat_68803;
    p55_concat_68954 <= p54_concat_68954;
    p55_concat_69913 <= p55_concat_69913_comb;
    p55_add_69216 <= p54_add_69216;
    p55_add_69255 <= p54_add_69255;
    p55_add_69945 <= p55_add_69945_comb;
  end

  // ===== Pipe stage 56:
  wire [31:0] p56_add_70003_comb;
  wire [31:0] p56_and_70008_comb;
  wire [31:0] p56_add_70004_comb;
  wire [31:0] p56_add_70005_comb;
  wire [31:0] p56_add_70027_comb;
  wire [31:0] p56_nor_70007_comb;
  wire [31:0] p56_add_70029_comb;
  wire [31:0] p56_add_70030_comb;
  assign p56_add_70003_comb = {p55_add_69880[5:0] ^ p55_add_69880[10:5] ^ p55_add_69880[24:19], p55_add_69880[31:27] ^ p55_add_69880[4:0] ^ p55_add_69880[18:14], p55_add_69880[26:13] ^ p55_add_69880[31:18] ^ p55_add_69880[13:0], p55_add_69880[12:6] ^ p55_add_69880[17:11] ^ p55_add_69880[31:25]} + (p55_add_69880 & p55_add_69793 ^ p55_nor_69882);
  assign p56_and_70008_comb = p55_add_69907 & p55_add_69816;
  assign p56_add_70004_comb = p56_add_70003_comb + p55_add_69885;
  assign p56_add_70005_comb = p56_add_70004_comb + p55_add_69729;
  assign p56_add_70027_comb = (p56_and_70008_comb ^ p55_add_69907 & p55_add_69729 ^ p55_and_69886) + p55_add_69879;
  assign p56_nor_70007_comb = ~(p56_add_70005_comb | ~p55_add_69793);
  assign p56_add_70029_comb = p56_add_70027_comb + {p55_add_69907[1:0] ^ p55_add_69907[12:11] ^ p55_add_69907[21:20], p55_add_69907[31:21] ^ p55_add_69907[10:0] ^ p55_add_69907[19:9], p55_add_69907[20:12] ^ p55_add_69907[31:23] ^ p55_add_69907[8:0], p55_add_69907[11:2] ^ p55_add_69907[22:13] ^ p55_add_69907[31:22]};
  assign p56_add_70030_comb = p55_concat_68803 + p55_add_69880;

  // Registers for pipe stage 56:
  reg [31:0] p56_add_67724;
  reg [31:0] p56_add_67758;
  reg [31:0] p56_add_69880;
  reg [31:0] p56_add_70004;
  reg [31:0] p56_add_70005;
  reg [31:0] p56_nor_70007;
  reg [31:0] p56_add_69813;
  reg [31:0] p56_add_69816;
  reg [31:0] p56_add_69907;
  reg [31:0] p56_add_69908;
  reg [31:0] p56_and_70008;
  reg [31:0] p56_add_70029;
  reg [31:0] p56_add_70030;
  reg [31:0] p56_concat_68954;
  reg [31:0] p56_concat_69913;
  reg [31:0] p56_add_69216;
  reg [31:0] p56_add_69255;
  reg [31:0] p56_add_69945;
  always_ff @ (posedge clk) begin
    p56_add_67724 <= p55_add_67724;
    p56_add_67758 <= p55_add_67758;
    p56_add_69880 <= p55_add_69880;
    p56_add_70004 <= p56_add_70004_comb;
    p56_add_70005 <= p56_add_70005_comb;
    p56_nor_70007 <= p56_nor_70007_comb;
    p56_add_69813 <= p55_add_69813;
    p56_add_69816 <= p55_add_69816;
    p56_add_69907 <= p55_add_69907;
    p56_add_69908 <= p55_add_69908;
    p56_and_70008 <= p56_and_70008_comb;
    p56_add_70029 <= p56_add_70029_comb;
    p56_add_70030 <= p56_add_70030_comb;
    p56_concat_68954 <= p55_concat_68954;
    p56_concat_69913 <= p55_concat_69913;
    p56_add_69216 <= p55_add_69216;
    p56_add_69255 <= p55_add_69255;
    p56_add_69945 <= p55_add_69945;
  end

  // ===== Pipe stage 57:
  wire [31:0] p57_add_70086_comb;
  wire [31:0] p57_and_70091_comb;
  wire [31:0] p57_add_70087_comb;
  wire [31:0] p57_add_70088_comb;
  wire [31:0] p57_add_70110_comb;
  wire [31:0] p57_nor_70090_comb;
  wire [31:0] p57_add_70112_comb;
  wire [31:0] p57_add_70113_comb;
  assign p57_add_70086_comb = (p56_add_70005 & p56_add_69880 ^ p56_nor_70007) + {p56_add_70005[5:0] ^ p56_add_70005[10:5] ^ p56_add_70005[24:19], p56_add_70005[31:27] ^ p56_add_70005[4:0] ^ p56_add_70005[18:14], p56_add_70005[26:13] ^ p56_add_70005[31:18] ^ p56_add_70005[13:0], p56_add_70005[12:6] ^ p56_add_70005[17:11] ^ p56_add_70005[31:25]};
  assign p57_and_70091_comb = p56_add_70029 & p56_add_69907;
  assign p57_add_70087_comb = p57_add_70086_comb + p56_add_69813;
  assign p57_add_70088_comb = p57_add_70087_comb + p56_add_69816;
  assign p57_add_70110_comb = (p57_and_70091_comb ^ p56_add_70029 & p56_add_69816 ^ p56_and_70008) + p56_add_70004;
  assign p57_nor_70090_comb = ~(p57_add_70088_comb | ~p56_add_69880);
  assign p57_add_70112_comb = p57_add_70110_comb + {p56_add_70029[1:0] ^ p56_add_70029[12:11] ^ p56_add_70029[21:20], p56_add_70029[31:21] ^ p56_add_70029[10:0] ^ p56_add_70029[19:9], p56_add_70029[20:12] ^ p56_add_70029[31:23] ^ p56_add_70029[8:0], p56_add_70029[11:2] ^ p56_add_70029[22:13] ^ p56_add_70029[31:22]};
  assign p57_add_70113_comb = p56_concat_68954 + p56_add_70005;

  // Registers for pipe stage 57:
  reg [31:0] p57_add_67724;
  reg [31:0] p57_add_67758;
  reg [31:0] p57_add_70005;
  reg [31:0] p57_add_70087;
  reg [31:0] p57_add_70088;
  reg [31:0] p57_nor_70090;
  reg [31:0] p57_add_69907;
  reg [31:0] p57_add_69908;
  reg [31:0] p57_add_70029;
  reg [31:0] p57_and_70091;
  reg [31:0] p57_add_70030;
  reg [31:0] p57_add_70112;
  reg [31:0] p57_add_70113;
  reg [31:0] p57_concat_69913;
  reg [31:0] p57_add_69216;
  reg [31:0] p57_add_69255;
  reg [31:0] p57_add_69945;
  always_ff @ (posedge clk) begin
    p57_add_67724 <= p56_add_67724;
    p57_add_67758 <= p56_add_67758;
    p57_add_70005 <= p56_add_70005;
    p57_add_70087 <= p57_add_70087_comb;
    p57_add_70088 <= p57_add_70088_comb;
    p57_nor_70090 <= p57_nor_70090_comb;
    p57_add_69907 <= p56_add_69907;
    p57_add_69908 <= p56_add_69908;
    p57_add_70029 <= p56_add_70029;
    p57_and_70091 <= p57_and_70091_comb;
    p57_add_70030 <= p56_add_70030;
    p57_add_70112 <= p57_add_70112_comb;
    p57_add_70113 <= p57_add_70113_comb;
    p57_concat_69913 <= p56_concat_69913;
    p57_add_69216 <= p56_add_69216;
    p57_add_69255 <= p56_add_69255;
    p57_add_69945 <= p56_add_69945;
  end

  // ===== Pipe stage 58:
  wire [31:0] p58_add_70167_comb;
  wire [31:0] p58_and_70172_comb;
  wire [31:0] p58_add_70168_comb;
  wire [31:0] p58_add_70169_comb;
  wire [31:0] p58_add_70191_comb;
  wire [31:0] p58_nor_70171_comb;
  wire [31:0] p58_add_70193_comb;
  wire [31:0] p58_add_70194_comb;
  assign p58_add_70167_comb = {p57_add_70088[5:0] ^ p57_add_70088[10:5] ^ p57_add_70088[24:19], p57_add_70088[31:27] ^ p57_add_70088[4:0] ^ p57_add_70088[18:14], p57_add_70088[26:13] ^ p57_add_70088[31:18] ^ p57_add_70088[13:0], p57_add_70088[12:6] ^ p57_add_70088[17:11] ^ p57_add_70088[31:25]} + (p57_add_70088 & p57_add_70005 ^ p57_nor_70090);
  assign p58_and_70172_comb = p57_add_70112 & p57_add_70029;
  assign p58_add_70168_comb = p58_add_70167_comb + p57_add_69908;
  assign p58_add_70169_comb = p58_add_70168_comb + p57_add_69907;
  assign p58_add_70191_comb = (p58_and_70172_comb ^ p57_add_70112 & p57_add_69907 ^ p57_and_70091) + p57_add_70087;
  assign p58_nor_70171_comb = ~(p58_add_70169_comb | ~p57_add_70005);
  assign p58_add_70193_comb = p58_add_70191_comb + {p57_add_70112[1:0] ^ p57_add_70112[12:11] ^ p57_add_70112[21:20], p57_add_70112[31:21] ^ p57_add_70112[10:0] ^ p57_add_70112[19:9], p57_add_70112[20:12] ^ p57_add_70112[31:23] ^ p57_add_70112[8:0], p57_add_70112[11:2] ^ p57_add_70112[22:13] ^ p57_add_70112[31:22]};
  assign p58_add_70194_comb = p57_concat_69913 + p57_add_70088;

  // Registers for pipe stage 58:
  reg [31:0] p58_add_67724;
  reg [31:0] p58_add_67758;
  reg [31:0] p58_add_70088;
  reg [31:0] p58_add_70168;
  reg [31:0] p58_add_70169;
  reg [31:0] p58_add_70029;
  reg [31:0] p58_nor_70171;
  reg [31:0] p58_add_70030;
  reg [31:0] p58_add_70112;
  reg [31:0] p58_and_70172;
  reg [31:0] p58_add_70193;
  reg [31:0] p58_add_70113;
  reg [31:0] p58_add_70194;
  reg [31:0] p58_add_69216;
  reg [31:0] p58_add_69255;
  reg [31:0] p58_add_69945;
  always_ff @ (posedge clk) begin
    p58_add_67724 <= p57_add_67724;
    p58_add_67758 <= p57_add_67758;
    p58_add_70088 <= p57_add_70088;
    p58_add_70168 <= p58_add_70168_comb;
    p58_add_70169 <= p58_add_70169_comb;
    p58_add_70029 <= p57_add_70029;
    p58_nor_70171 <= p58_nor_70171_comb;
    p58_add_70030 <= p57_add_70030;
    p58_add_70112 <= p57_add_70112;
    p58_and_70172 <= p58_and_70172_comb;
    p58_add_70193 <= p58_add_70193_comb;
    p58_add_70113 <= p57_add_70113;
    p58_add_70194 <= p58_add_70194_comb;
    p58_add_69216 <= p57_add_69216;
    p58_add_69255 <= p57_add_69255;
    p58_add_69945 <= p57_add_69945;
  end

  // ===== Pipe stage 59:
  wire [31:0] p59_add_70246_comb;
  wire [31:0] p59_and_70251_comb;
  wire [31:0] p59_add_70247_comb;
  wire [31:0] p59_add_70248_comb;
  wire [31:0] p59_add_70270_comb;
  wire [31:0] p59_nor_70250_comb;
  wire [31:0] p59_add_70272_comb;
  wire [31:0] p59_add_70273_comb;
  assign p59_add_70246_comb = (p58_add_70169 & p58_add_70088 ^ p58_nor_70171) + {p58_add_70169[5:0] ^ p58_add_70169[10:5] ^ p58_add_70169[24:19], p58_add_70169[31:27] ^ p58_add_70169[4:0] ^ p58_add_70169[18:14], p58_add_70169[26:13] ^ p58_add_70169[31:18] ^ p58_add_70169[13:0], p58_add_70169[12:6] ^ p58_add_70169[17:11] ^ p58_add_70169[31:25]};
  assign p59_and_70251_comb = p58_add_70193 & p58_add_70112;
  assign p59_add_70247_comb = p59_add_70246_comb + p58_add_70030;
  assign p59_add_70248_comb = p59_add_70247_comb + p58_add_70029;
  assign p59_add_70270_comb = (p59_and_70251_comb ^ p58_add_70193 & p58_add_70029 ^ p58_and_70172) + p58_add_70168;
  assign p59_nor_70250_comb = ~(p59_add_70248_comb | ~p58_add_70088);
  assign p59_add_70272_comb = p59_add_70270_comb + {p58_add_70193[1:0] ^ p58_add_70193[12:11] ^ p58_add_70193[21:20], p58_add_70193[31:21] ^ p58_add_70193[10:0] ^ p58_add_70193[19:9], p58_add_70193[20:12] ^ p58_add_70193[31:23] ^ p58_add_70193[8:0], p58_add_70193[11:2] ^ p58_add_70193[22:13] ^ p58_add_70193[31:22]};
  assign p59_add_70273_comb = p58_add_70169 + p58_add_69216;

  // Registers for pipe stage 59:
  reg [31:0] p59_add_67724;
  reg [31:0] p59_add_67758;
  reg [31:0] p59_add_70169;
  reg [31:0] p59_add_70247;
  reg [31:0] p59_add_70112;
  reg [31:0] p59_add_70248;
  reg [31:0] p59_nor_70250;
  reg [31:0] p59_add_70193;
  reg [31:0] p59_add_70113;
  reg [31:0] p59_and_70251;
  reg [31:0] p59_add_70272;
  reg [31:0] p59_add_70194;
  reg [31:0] p59_add_70273;
  reg [31:0] p59_add_69255;
  reg [31:0] p59_add_69945;
  always_ff @ (posedge clk) begin
    p59_add_67724 <= p58_add_67724;
    p59_add_67758 <= p58_add_67758;
    p59_add_70169 <= p58_add_70169;
    p59_add_70247 <= p59_add_70247_comb;
    p59_add_70112 <= p58_add_70112;
    p59_add_70248 <= p59_add_70248_comb;
    p59_nor_70250 <= p59_nor_70250_comb;
    p59_add_70193 <= p58_add_70193;
    p59_add_70113 <= p58_add_70113;
    p59_and_70251 <= p59_and_70251_comb;
    p59_add_70272 <= p59_add_70272_comb;
    p59_add_70194 <= p58_add_70194;
    p59_add_70273 <= p59_add_70273_comb;
    p59_add_69255 <= p58_add_69255;
    p59_add_69945 <= p58_add_69945;
  end

  // ===== Pipe stage 60:
  wire [31:0] p60_add_70323_comb;
  wire [31:0] p60_and_70328_comb;
  wire [31:0] p60_add_70324_comb;
  wire [31:0] p60_add_70325_comb;
  wire [31:0] p60_add_70347_comb;
  wire [31:0] p60_nor_70327_comb;
  wire [31:0] p60_add_70349_comb;
  wire [31:0] p60_add_70350_comb;
  assign p60_add_70323_comb = (p59_add_70248 & p59_add_70169 ^ p59_nor_70250) + {p59_add_70248[5:0] ^ p59_add_70248[10:5] ^ p59_add_70248[24:19], p59_add_70248[31:27] ^ p59_add_70248[4:0] ^ p59_add_70248[18:14], p59_add_70248[26:13] ^ p59_add_70248[31:18] ^ p59_add_70248[13:0], p59_add_70248[12:6] ^ p59_add_70248[17:11] ^ p59_add_70248[31:25]};
  assign p60_and_70328_comb = p59_add_70272 & p59_add_70193;
  assign p60_add_70324_comb = p60_add_70323_comb + p59_add_70113;
  assign p60_add_70325_comb = p60_add_70324_comb + p59_add_70112;
  assign p60_add_70347_comb = (p60_and_70328_comb ^ p59_add_70272 & p59_add_70112 ^ p59_and_70251) + p59_add_70247;
  assign p60_nor_70327_comb = ~(p60_add_70325_comb | ~p59_add_70169);
  assign p60_add_70349_comb = p60_add_70347_comb + {p59_add_70272[1:0] ^ p59_add_70272[12:11] ^ p59_add_70272[21:20], p59_add_70272[31:21] ^ p59_add_70272[10:0] ^ p59_add_70272[19:9], p59_add_70272[20:12] ^ p59_add_70272[31:23] ^ p59_add_70272[8:0], p59_add_70272[11:2] ^ p59_add_70272[22:13] ^ p59_add_70272[31:22]};
  assign p60_add_70350_comb = p59_add_67724 + p59_add_70248;

  // Registers for pipe stage 60:
  reg [31:0] p60_add_67758;
  reg [31:0] p60_add_70248;
  reg [31:0] p60_add_70193;
  reg [31:0] p60_add_70324;
  reg [31:0] p60_add_70325;
  reg [31:0] p60_add_70272;
  reg [31:0] p60_nor_70327;
  reg [31:0] p60_and_70328;
  reg [31:0] p60_add_70194;
  reg [31:0] p60_add_70349;
  reg [31:0] p60_add_70273;
  reg [31:0] p60_add_69255;
  reg [31:0] p60_add_70350;
  reg [31:0] p60_add_69945;
  always_ff @ (posedge clk) begin
    p60_add_67758 <= p59_add_67758;
    p60_add_70248 <= p59_add_70248;
    p60_add_70193 <= p59_add_70193;
    p60_add_70324 <= p60_add_70324_comb;
    p60_add_70325 <= p60_add_70325_comb;
    p60_add_70272 <= p59_add_70272;
    p60_nor_70327 <= p60_nor_70327_comb;
    p60_and_70328 <= p60_and_70328_comb;
    p60_add_70194 <= p59_add_70194;
    p60_add_70349 <= p60_add_70349_comb;
    p60_add_70273 <= p59_add_70273;
    p60_add_69255 <= p59_add_69255;
    p60_add_70350 <= p60_add_70350_comb;
    p60_add_69945 <= p59_add_69945;
  end

  // ===== Pipe stage 61:
  wire [31:0] p61_add_70398_comb;
  wire [31:0] p61_and_70401_comb;
  wire [31:0] p61_add_70399_comb;
  wire [31:0] p61_add_70400_comb;
  wire [31:0] p61_add_70422_comb;
  wire [31:0] p61_nor_70421_comb;
  wire [31:0] p61_add_70424_comb;
  wire [31:0] p61_add_70425_comb;
  assign p61_add_70398_comb = (p60_add_70325 & p60_add_70248 ^ p60_nor_70327) + {p60_add_70325[5:0] ^ p60_add_70325[10:5] ^ p60_add_70325[24:19], p60_add_70325[31:27] ^ p60_add_70325[4:0] ^ p60_add_70325[18:14], p60_add_70325[26:13] ^ p60_add_70325[31:18] ^ p60_add_70325[13:0], p60_add_70325[12:6] ^ p60_add_70325[17:11] ^ p60_add_70325[31:25]};
  assign p61_and_70401_comb = p60_add_70349 & p60_add_70272;
  assign p61_add_70399_comb = p61_add_70398_comb + p60_add_70194;
  assign p61_add_70400_comb = p61_add_70399_comb + p60_add_70193;
  assign p61_add_70422_comb = (p61_and_70401_comb ^ p60_add_70349 & p60_add_70193 ^ p60_and_70328) + p60_add_70324;
  assign p61_nor_70421_comb = ~(p61_add_70400_comb | ~p60_add_70248);
  assign p61_add_70424_comb = p61_add_70422_comb + {p60_add_70349[1:0] ^ p60_add_70349[12:11] ^ p60_add_70349[21:20], p60_add_70349[31:21] ^ p60_add_70349[10:0] ^ p60_add_70349[19:9], p60_add_70349[20:12] ^ p60_add_70349[31:23] ^ p60_add_70349[8:0], p60_add_70349[11:2] ^ p60_add_70349[22:13] ^ p60_add_70349[31:22]};
  assign p61_add_70425_comb = p60_add_67758 + p60_add_70325;

  // Registers for pipe stage 61:
  reg [31:0] p61_add_70325;
  reg [31:0] p61_add_70272;
  reg [31:0] p61_add_70399;
  reg [31:0] p61_add_70349;
  reg [31:0] p61_add_70400;
  reg [31:0] p61_and_70401;
  reg [31:0] p61_nor_70421;
  reg [31:0] p61_add_70424;
  reg [31:0] p61_add_70273;
  reg [31:0] p61_add_70425;
  reg [31:0] p61_add_69255;
  reg [31:0] p61_add_70350;
  reg [31:0] p61_add_69945;
  always_ff @ (posedge clk) begin
    p61_add_70325 <= p60_add_70325;
    p61_add_70272 <= p60_add_70272;
    p61_add_70399 <= p61_add_70399_comb;
    p61_add_70349 <= p60_add_70349;
    p61_add_70400 <= p61_add_70400_comb;
    p61_and_70401 <= p61_and_70401_comb;
    p61_nor_70421 <= p61_nor_70421_comb;
    p61_add_70424 <= p61_add_70424_comb;
    p61_add_70273 <= p60_add_70273;
    p61_add_70425 <= p61_add_70425_comb;
    p61_add_69255 <= p60_add_69255;
    p61_add_70350 <= p60_add_70350;
    p61_add_69945 <= p60_add_69945;
  end

  // ===== Pipe stage 62:
  wire [31:0] p62_and_70472_comb;
  wire [31:0] p62_add_70471_comb;
  wire [31:0] p62_add_70486_comb;
  wire [31:0] p62_add_70493_comb;
  wire [31:0] p62_add_70492_comb;
  wire [31:0] p62_add_70496_comb;
  wire [31:0] p62_nor_70497_comb;
  assign p62_and_70472_comb = p61_add_70424 & p61_add_70349;
  assign p62_add_70471_comb = {p61_add_70400[5:0] ^ p61_add_70400[10:5] ^ p61_add_70400[24:19], p61_add_70400[31:27] ^ p61_add_70400[4:0] ^ p61_add_70400[18:14], p61_add_70400[26:13] ^ p61_add_70400[31:18] ^ p61_add_70400[13:0], p61_add_70400[12:6] ^ p61_add_70400[17:11] ^ p61_add_70400[31:25]} + (p61_add_70400 & p61_add_70325 ^ p61_nor_70421);
  assign p62_add_70486_comb = p62_add_70471_comb + p61_add_70273;
  assign p62_add_70493_comb = (p62_and_70472_comb ^ p61_add_70424 & p61_add_70272 ^ p61_and_70401) + p61_add_70399;
  assign p62_add_70492_comb = p62_add_70486_comb + p61_add_70272;
  assign p62_add_70496_comb = p62_add_70493_comb + {p61_add_70424[1:0] ^ p61_add_70424[12:11] ^ p61_add_70424[21:20], p61_add_70424[31:21] ^ p61_add_70424[10:0] ^ p61_add_70424[19:9], p61_add_70424[20:12] ^ p61_add_70424[31:23] ^ p61_add_70424[8:0], p61_add_70424[11:2] ^ p61_add_70424[22:13] ^ p61_add_70424[31:22]};
  assign p62_nor_70497_comb = ~(p62_add_70492_comb | ~p61_add_70325);

  // Registers for pipe stage 62:
  reg [31:0] p62_add_70349;
  reg [31:0] p62_add_70400;
  reg [31:0] p62_add_70424;
  reg [31:0] p62_and_70472;
  reg [31:0] p62_add_70486;
  reg [31:0] p62_add_70492;
  reg [31:0] p62_add_70496;
  reg [31:0] p62_nor_70497;
  reg [31:0] p62_add_70425;
  reg [31:0] p62_add_69255;
  reg [31:0] p62_add_70350;
  reg [31:0] p62_add_69945;
  always_ff @ (posedge clk) begin
    p62_add_70349 <= p61_add_70349;
    p62_add_70400 <= p61_add_70400;
    p62_add_70424 <= p61_add_70424;
    p62_and_70472 <= p62_and_70472_comb;
    p62_add_70486 <= p62_add_70486_comb;
    p62_add_70492 <= p62_add_70492_comb;
    p62_add_70496 <= p62_add_70496_comb;
    p62_nor_70497 <= p62_nor_70497_comb;
    p62_add_70425 <= p61_add_70425;
    p62_add_69255 <= p61_add_69255;
    p62_add_70350 <= p61_add_70350;
    p62_add_69945 <= p61_add_69945;
  end

  // ===== Pipe stage 63:
  wire [31:0] p63_and_70539_comb;
  wire [31:0] p63_add_70560_comb;
  wire [31:0] p63_add_70561_comb;
  wire [31:0] p63_add_70563_comb;
  wire [31:0] p63_add_70564_comb;
  wire [31:0] p63_add_70565_comb;
  assign p63_and_70539_comb = p62_add_70496 & p62_add_70424;
  assign p63_add_70560_comb = {p62_add_70492[5:0] ^ p62_add_70492[10:5] ^ p62_add_70492[24:19], p62_add_70492[31:27] ^ p62_add_70492[4:0] ^ p62_add_70492[18:14], p62_add_70492[26:13] ^ p62_add_70492[31:18] ^ p62_add_70492[13:0], p62_add_70492[12:6] ^ p62_add_70492[17:11] ^ p62_add_70492[31:25]} + (p62_add_70492 & p62_add_70400 ^ p62_nor_70497);
  assign p63_add_70561_comb = (p63_and_70539_comb ^ p62_add_70496 & p62_add_70349 ^ p62_and_70472) + p62_add_70486;
  assign p63_add_70563_comb = p62_add_70350 + p63_add_70560_comb;
  assign p63_add_70564_comb = p63_add_70561_comb + {p62_add_70496[1:0] ^ p62_add_70496[12:11] ^ p62_add_70496[21:20], p62_add_70496[31:21] ^ p62_add_70496[10:0] ^ p62_add_70496[19:9], p62_add_70496[20:12] ^ p62_add_70496[31:23] ^ p62_add_70496[8:0], p62_add_70496[11:2] ^ p62_add_70496[22:13] ^ p62_add_70496[31:22]};
  assign p63_add_70565_comb = p63_add_70563_comb + p62_add_69945;

  // Registers for pipe stage 63:
  reg [31:0] p63_add_70349;
  reg [31:0] p63_add_70400;
  reg [31:0] p63_add_70424;
  reg [31:0] p63_add_70492;
  reg [31:0] p63_add_70496;
  reg [31:0] p63_and_70539;
  reg [31:0] p63_add_70564;
  reg [31:0] p63_add_70425;
  reg [31:0] p63_add_69255;
  reg [31:0] p63_add_70565;
  always_ff @ (posedge clk) begin
    p63_add_70349 <= p62_add_70349;
    p63_add_70400 <= p62_add_70400;
    p63_add_70424 <= p62_add_70424;
    p63_add_70492 <= p62_add_70492;
    p63_add_70496 <= p62_add_70496;
    p63_and_70539 <= p63_and_70539_comb;
    p63_add_70564 <= p63_add_70564_comb;
    p63_add_70425 <= p62_add_70425;
    p63_add_69255 <= p62_add_69255;
    p63_add_70565 <= p63_add_70565_comb;
  end

  // ===== Pipe stage 64:
  wire [31:0] p64_and_70586_comb;
  wire [31:0] p64_add_70600_comb;
  wire [31:0] p64_add_70619_comb;
  wire [31:0] p64_add_70627_comb;
  wire [30:0] p64_add_70641_comb;
  wire [30:0] p64_add_70643_comb;
  wire [29:0] p64_add_70645_comb;
  wire [31:0] p64_add_70630_comb;
  wire [31:0] p64_xor_70634_comb;
  wire [31:0] p64_concat_70649_comb;
  wire [31:0] p64_concat_70650_comb;
  wire [31:0] p64_concat_70651_comb;
  wire [31:0] p64_add_70652_comb;
  wire [31:0] p64_add_70653_comb;
  wire [31:0] p64_add_70633_comb;
  assign p64_and_70586_comb = p63_add_70564 & p63_add_70496;
  assign p64_add_70600_comb = p63_add_70565 + p63_add_70349;
  assign p64_add_70619_comb = (p64_and_70586_comb ^ p63_add_70564 & p63_add_70424 ^ p63_and_70539) + p63_add_70565;
  assign p64_add_70627_comb = p64_add_70619_comb + {p63_add_70564[1:0] ^ p63_add_70564[12:11] ^ p63_add_70564[21:20], p63_add_70564[31:21] ^ p63_add_70564[10:0] ^ p63_add_70564[19:9], p63_add_70564[20:12] ^ p63_add_70564[31:23] ^ p63_add_70564[8:0], p63_add_70564[11:2] ^ p63_add_70564[22:13] ^ p63_add_70564[31:22]};
  assign p64_add_70641_comb = p63_add_70564[31:1] + 31'h1e37_79b9;
  assign p64_add_70643_comb = p63_add_70496[31:1] + 31'h52a7_fa9d;
  assign p64_add_70645_comb = p64_add_70600_comb[31:2] + 30'h26c1_5a23;
  assign p64_add_70630_comb = {p64_add_70600_comb[5:0] ^ p64_add_70600_comb[10:5] ^ p64_add_70600_comb[24:19], p64_add_70600_comb[31:27] ^ p64_add_70600_comb[4:0] ^ p64_add_70600_comb[18:14], p64_add_70600_comb[26:13] ^ p64_add_70600_comb[31:18] ^ p64_add_70600_comb[13:0], p64_add_70600_comb[12:6] ^ p64_add_70600_comb[17:11] ^ p64_add_70600_comb[31:25]} + (p64_add_70600_comb & p63_add_70492 ^ ~(p64_add_70600_comb | ~p63_add_70400));
  assign p64_xor_70634_comb = p64_add_70627_comb & p63_add_70564 ^ p64_add_70627_comb & p63_add_70496 ^ p64_and_70586_comb;
  assign p64_concat_70649_comb = {p64_add_70641_comb, p63_add_70564[0]};
  assign p64_concat_70650_comb = {p64_add_70643_comb, p63_add_70496[0]};
  assign p64_concat_70651_comb = {p64_add_70645_comb, p64_add_70600_comb[1:0]};
  assign p64_add_70652_comb = p63_add_70492 + 32'h1f83_d9ab;
  assign p64_add_70653_comb = p63_add_70400 + 32'h5be0_cd19;
  assign p64_add_70633_comb = p63_add_70425 + p64_add_70630_comb;

  // Registers for pipe stage 64:
  reg [31:0] p64_add_70424;
  reg [31:0] p64_add_70627;
  reg [31:0] p64_xor_70634;
  reg [31:0] p64_concat_70649;
  reg [31:0] p64_concat_70650;
  reg [31:0] p64_concat_70651;
  reg [31:0] p64_add_70652;
  reg [31:0] p64_add_70653;
  reg [31:0] p64_add_70633;
  reg [31:0] p64_add_69255;
  always_ff @ (posedge clk) begin
    p64_add_70424 <= p63_add_70424;
    p64_add_70627 <= p64_add_70627_comb;
    p64_xor_70634 <= p64_xor_70634_comb;
    p64_concat_70649 <= p64_concat_70649_comb;
    p64_concat_70650 <= p64_concat_70650_comb;
    p64_concat_70651 <= p64_concat_70651_comb;
    p64_add_70652 <= p64_add_70652_comb;
    p64_add_70653 <= p64_add_70653_comb;
    p64_add_70633 <= p64_add_70633_comb;
    p64_add_69255 <= p63_add_69255;
  end

  // ===== Pipe stage 65:
  wire [31:0] p65_add_70691_comb;
  wire [31:0] p65_add_70694_comb;
  wire [31:0] p65_add_70695_comb;
  wire [31:0] p65_add_70697_comb;
  wire [31:0] p65_add_70698_comb;
  wire [31:0] p65_add_70699_comb;
  wire [31:0] p65_add_70700_comb;
  wire [255:0] p65_tuple_70701_comb;
  assign p65_add_70691_comb = p64_add_70633 + p64_add_69255;
  assign p65_add_70694_comb = p64_xor_70634 + {p64_add_70627[1:0] ^ p64_add_70627[12:11] ^ p64_add_70627[21:20], p64_add_70627[31:21] ^ p64_add_70627[10:0] ^ p64_add_70627[19:9], p64_add_70627[20:12] ^ p64_add_70627[31:23] ^ p64_add_70627[8:0], p64_add_70627[11:2] ^ p64_add_70627[22:13] ^ p64_add_70627[31:22]};
  assign p65_add_70695_comb = p65_add_70691_comb + 32'h6a09_e667;
  assign p65_add_70697_comb = p65_add_70691_comb + 32'h510e_527f;
  assign p65_add_70698_comb = p65_add_70694_comb + p65_add_70695_comb;
  assign p65_add_70699_comb = p64_add_70627 + 32'hbb67_ae85;
  assign p65_add_70700_comb = p65_add_70697_comb + p64_add_70424;
  assign p65_tuple_70701_comb = {p65_add_70698_comb, p65_add_70699_comb, p64_concat_70649, p64_concat_70650, p65_add_70700_comb, p64_concat_70651, p64_add_70652, p64_add_70653};

  // Registers for pipe stage 65:
  reg [255:0] p65_tuple_70701;
  always_ff @ (posedge clk) begin
    p65_tuple_70701 <= p65_tuple_70701_comb;
  end
  assign out = p65_tuple_70701;
endmodule
