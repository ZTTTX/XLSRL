module xls_test(
  input wire clk,
  input wire [511:0] message,
  output wire [255:0] out
);
  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [511:0] p0_message;
  always_ff @ (posedge clk) begin
    p0_message <= message;
  end

  // ===== Pipe stage 1:
  wire [28:0] p1_add_63010_comb;
  wire [30:0] p1_add_63014_comb;
  wire p1_bit_slice_63016_comb;
  wire [31:0] p1_concat_63033_comb;
  wire [29:0] p1_add_63040_comb;
  wire [31:0] p1_xor_63046_comb;
  wire [31:0] p1_add_63047_comb;
  assign p1_add_63010_comb = p0_message[511:483] + 29'h1e6e_fdad;
  assign p1_add_63014_comb = {p1_add_63010_comb, p0_message[482:481]} + 31'h52a7_fa9d;
  assign p1_bit_slice_63016_comb = p0_message[480];
  assign p1_concat_63033_comb = {p1_add_63014_comb, p1_bit_slice_63016_comb};
  assign p1_add_63040_comb = p0_message[479:450] + 30'h242e_c78f;
  assign p1_xor_63046_comb = p1_concat_63033_comb & 32'h510e_527f ^ ~(p1_concat_63033_comb | 32'h64fa_9773);
  assign p1_add_63047_comb = {{p1_add_63014_comb[4:0], p1_bit_slice_63016_comb} ^ p1_add_63014_comb[9:4] ^ p1_add_63014_comb[23:18], p1_add_63014_comb[30:26] ^ {p1_add_63014_comb[3:0], p1_bit_slice_63016_comb} ^ p1_add_63014_comb[17:13], p1_add_63014_comb[25:12] ^ p1_add_63014_comb[30:17] ^ {p1_add_63014_comb[12:0], p1_bit_slice_63016_comb}, p1_add_63014_comb[11:5] ^ p1_add_63014_comb[16:10] ^ p1_add_63014_comb[30:24]} + {p1_add_63040_comb, p0_message[449:448]};

  // Registers for pipe stage 1:
  reg [511:0] p1_message;
  reg [28:0] p1_add_63010;
  reg [30:0] p1_add_63014;
  reg p1_bit_slice_63016;
  reg [31:0] p1_concat_63033;
  reg [31:0] p1_xor_63046;
  reg [31:0] p1_add_63047;
  always_ff @ (posedge clk) begin
    p1_message <= p0_message;
    p1_add_63010 <= p1_add_63010_comb;
    p1_add_63014 <= p1_add_63014_comb;
    p1_bit_slice_63016 <= p1_bit_slice_63016_comb;
    p1_concat_63033 <= p1_concat_63033_comb;
    p1_xor_63046 <= p1_xor_63046_comb;
    p1_add_63047 <= p1_add_63047_comb;
  end

  // ===== Pipe stage 2:
  wire [31:0] p2_add_63062_comb;
  wire [30:0] p2_add_63065_comb;
  wire [31:0] p2_concat_63072_comb;
  wire [31:0] p2_concat_63100_comb;
  wire [31:0] p2_concat_63103_comb;
  wire [31:0] p2_add_63120_comb;
  wire [31:0] p2_add_63096_comb;
  wire [31:0] p2_add_63097_comb;
  assign p2_add_63062_comb = p1_xor_63046 + p1_add_63047;
  assign p2_add_63065_comb = p2_add_63062_comb[31:1] + 31'h1e37_79b9;
  assign p2_concat_63072_comb = {p2_add_63065_comb, p2_add_63062_comb[0]};
  assign p2_concat_63100_comb = {~p1_add_63014, ~p1_bit_slice_63016};
  assign p2_concat_63103_comb = {~p2_add_63065_comb, ~p2_add_63062_comb[0]};
  assign p2_add_63120_comb = {p1_message[390:388] ^ p1_message[401:399], p1_message[387:384] ^ p1_message[398:395] ^ p1_message[415:412], p1_message[415:405] ^ p1_message[394:384] ^ p1_message[411:401], p1_message[404:391] ^ p1_message[415:402] ^ p1_message[400:387]} + p1_message[447:416];
  assign p2_add_63096_comb = ({p2_add_63065_comb & p1_add_63014, p2_add_63062_comb[0] & p1_bit_slice_63016} ^ ~(p2_concat_63072_comb | 32'haef1_ad80)) + {{p2_add_63065_comb[4:0], p2_add_63062_comb[0]} ^ p2_add_63065_comb[9:4] ^ p2_add_63065_comb[23:18], p2_add_63065_comb[30:26] ^ {p2_add_63065_comb[3:0], p2_add_63062_comb[0]} ^ p2_add_63065_comb[17:13], p2_add_63065_comb[25:12] ^ p2_add_63065_comb[30:17] ^ {p2_add_63065_comb[12:0], p2_add_63062_comb[0]}, p2_add_63065_comb[11:5] ^ p2_add_63065_comb[16:10] ^ p2_add_63065_comb[30:24]};
  assign p2_add_63097_comb = p1_message[447:416] + 32'h50c6_645b;

  // Registers for pipe stage 2:
  reg [511:0] p2_message;
  reg [28:0] p2_add_63010;
  reg [31:0] p2_concat_63033;
  reg [31:0] p2_add_63062;
  reg [31:0] p2_concat_63072;
  reg [31:0] p2_concat_63100;
  reg [31:0] p2_concat_63103;
  reg [31:0] p2_add_63120;
  reg [31:0] p2_add_63096;
  reg [31:0] p2_add_63097;
  always_ff @ (posedge clk) begin
    p2_message <= p1_message;
    p2_add_63010 <= p1_add_63010;
    p2_concat_63033 <= p1_concat_63033;
    p2_add_63062 <= p2_add_63062_comb;
    p2_concat_63072 <= p2_concat_63072_comb;
    p2_concat_63100 <= p2_concat_63100_comb;
    p2_concat_63103 <= p2_concat_63103_comb;
    p2_add_63120 <= p2_add_63120_comb;
    p2_add_63096 <= p2_add_63096_comb;
    p2_add_63097 <= p2_add_63097_comb;
  end

  // ===== Pipe stage 3:
  wire [31:0] p3_add_63141_comb;
  wire [31:0] p3_add_63143_comb;
  wire [29:0] p3_add_63162_comb;
  wire [31:0] p3_xor_63168_comb;
  wire [31:0] p3_add_63169_comb;
  assign p3_add_63141_comb = p2_add_63096 + p2_add_63097;
  assign p3_add_63143_comb = p3_add_63141_comb + 32'hbb67_ae85;
  assign p3_add_63162_comb = p2_message[415:386] + 30'h0eb1_0b89;
  assign p3_xor_63168_comb = p3_add_63143_comb & p2_concat_63072 ^ ~(p3_add_63143_comb | p2_concat_63100);
  assign p3_add_63169_comb = {p3_add_63143_comb[5:0] ^ p3_add_63143_comb[10:5] ^ p3_add_63143_comb[24:19], p3_add_63143_comb[31:27] ^ p3_add_63143_comb[4:0] ^ p3_add_63143_comb[18:14], p3_add_63143_comb[26:13] ^ p3_add_63143_comb[31:18] ^ p3_add_63143_comb[13:0], p3_add_63143_comb[12:6] ^ p3_add_63143_comb[17:11] ^ p3_add_63143_comb[31:25]} + {p3_add_63162_comb, p2_message[385:384]};

  // Registers for pipe stage 3:
  reg [511:0] p3_message;
  reg [28:0] p3_add_63010;
  reg [31:0] p3_concat_63033;
  reg [31:0] p3_add_63062;
  reg [31:0] p3_concat_63072;
  reg [31:0] p3_add_63143;
  reg [31:0] p3_xor_63168;
  reg [31:0] p3_add_63169;
  reg [31:0] p3_concat_63103;
  reg [31:0] p3_add_63120;
  reg [31:0] p3_add_63141;
  always_ff @ (posedge clk) begin
    p3_message <= p2_message;
    p3_add_63010 <= p2_add_63010;
    p3_concat_63033 <= p2_concat_63033;
    p3_add_63062 <= p2_add_63062;
    p3_concat_63072 <= p2_concat_63072;
    p3_add_63143 <= p3_add_63143_comb;
    p3_xor_63168 <= p3_xor_63168_comb;
    p3_add_63169 <= p3_add_63169_comb;
    p3_concat_63103 <= p2_concat_63103;
    p3_add_63120 <= p2_add_63120;
    p3_add_63141 <= p3_add_63141_comb;
  end

  // ===== Pipe stage 4:
  wire [31:0] p4_add_63192_comb;
  wire [31:0] p4_add_63219_comb;
  wire [31:0] p4_add_63194_comb;
  wire [31:0] p4_and_63238_comb;
  wire [31:0] p4_add_63243_comb;
  wire [31:0] p4_add_63216_comb;
  wire [31:0] p4_add_63244_comb;
  assign p4_add_63192_comb = p3_xor_63168 + p3_add_63169;
  assign p4_add_63219_comb = {p3_add_63010, p3_message[482:480]} + 32'h0890_9ae5;
  assign p4_add_63194_comb = p4_add_63192_comb + 32'h6a09_e667;
  assign p4_and_63238_comb = p4_add_63219_comb & 32'h6a09_e667;
  assign p4_add_63243_comb = {p4_add_63219_comb[1:0] ^ p4_add_63219_comb[12:11] ^ p4_add_63219_comb[21:20], p4_add_63219_comb[31:21] ^ p4_add_63219_comb[10:0] ^ p4_add_63219_comb[19:9], p4_add_63219_comb[20:12] ^ p4_add_63219_comb[31:23] ^ p4_add_63219_comb[8:0], p4_add_63219_comb[11:2] ^ p4_add_63219_comb[22:13] ^ p4_add_63219_comb[31:22]} + (p4_and_63238_comb ^ p4_add_63219_comb & 32'hbb67_ae85 ^ 32'h2a01_a605);
  assign p4_add_63216_comb = {p4_add_63194_comb[5:0] ^ p4_add_63194_comb[10:5] ^ p4_add_63194_comb[24:19], p4_add_63194_comb[31:27] ^ p4_add_63194_comb[4:0] ^ p4_add_63194_comb[18:14], p4_add_63194_comb[26:13] ^ p4_add_63194_comb[31:18] ^ p4_add_63194_comb[13:0], p4_add_63194_comb[12:6] ^ p4_add_63194_comb[17:11] ^ p4_add_63194_comb[31:25]} + (p4_add_63194_comb & p3_add_63143 ^ ~(p4_add_63194_comb | p3_concat_63103));
  assign p4_add_63244_comb = p3_add_63062 + p4_add_63243_comb;

  // Registers for pipe stage 4:
  reg [511:0] p4_message;
  reg [31:0] p4_concat_63033;
  reg [31:0] p4_concat_63072;
  reg [31:0] p4_add_63143;
  reg [31:0] p4_add_63192;
  reg [31:0] p4_add_63194;
  reg [31:0] p4_add_63216;
  reg [31:0] p4_add_63219;
  reg [31:0] p4_and_63238;
  reg [31:0] p4_add_63244;
  reg [31:0] p4_add_63120;
  reg [31:0] p4_add_63141;
  always_ff @ (posedge clk) begin
    p4_message <= p3_message;
    p4_concat_63033 <= p3_concat_63033;
    p4_concat_63072 <= p3_concat_63072;
    p4_add_63143 <= p3_add_63143;
    p4_add_63192 <= p4_add_63192_comb;
    p4_add_63194 <= p4_add_63194_comb;
    p4_add_63216 <= p4_add_63216_comb;
    p4_add_63219 <= p4_add_63219_comb;
    p4_and_63238 <= p4_and_63238_comb;
    p4_add_63244 <= p4_add_63244_comb;
    p4_add_63120 <= p3_add_63120;
    p4_add_63141 <= p3_add_63141;
  end

  // ===== Pipe stage 5:
  wire [31:0] p5_and_63292_comb;
  wire [31:0] p5_add_63296_comb;
  wire [31:0] p5_add_63271_comb;
  wire [31:0] p5_add_63272_comb;
  wire [31:0] p5_add_63297_comb;
  wire [31:0] p5_add_63273_comb;
  wire [31:0] p5_and_63298_comb;
  wire [31:0] p5_add_63274_comb;
  wire [31:0] p5_xor_63300_comb;
  wire [31:0] p5_add_63317_comb;
  assign p5_and_63292_comb = p4_add_63244 & p4_add_63219;
  assign p5_add_63296_comb = {p4_add_63244[1:0] ^ p4_add_63244[12:11] ^ p4_add_63244[21:20], p4_add_63244[31:21] ^ p4_add_63244[10:0] ^ p4_add_63244[19:9], p4_add_63244[20:12] ^ p4_add_63244[31:23] ^ p4_add_63244[8:0], p4_add_63244[11:2] ^ p4_add_63244[22:13] ^ p4_add_63244[31:22]} + (p5_and_63292_comb ^ p4_add_63244 & 32'h6a09_e667 ^ p4_and_63238);
  assign p5_add_63271_comb = p4_add_63216 + 32'h3956_c25b;
  assign p5_add_63272_comb = p4_concat_63033 + p4_message[383:352];
  assign p5_add_63297_comb = p4_add_63141 + p5_add_63296_comb;
  assign p5_add_63273_comb = p5_add_63271_comb + p5_add_63272_comb;
  assign p5_and_63298_comb = p5_add_63297_comb & p4_add_63244;
  assign p5_add_63274_comb = p4_add_63219 + p5_add_63273_comb;
  assign p5_xor_63300_comb = p5_and_63298_comb ^ p5_add_63297_comb & p4_add_63219 ^ p5_and_63292_comb;
  assign p5_add_63317_comb = {p4_message[326:324] ^ p4_message[337:335], p4_message[323:320] ^ p4_message[334:331] ^ p4_message[351:348], p4_message[351:341] ^ p4_message[330:320] ^ p4_message[347:337], p4_message[340:327] ^ p4_message[351:338] ^ p4_message[336:323]} + p4_message[383:352];

  // Registers for pipe stage 5:
  reg [511:0] p5_message;
  reg [31:0] p5_concat_63072;
  reg [31:0] p5_add_63143;
  reg [31:0] p5_add_63192;
  reg [31:0] p5_add_63194;
  reg [31:0] p5_add_63273;
  reg [31:0] p5_add_63274;
  reg [31:0] p5_add_63244;
  reg [31:0] p5_add_63297;
  reg [31:0] p5_and_63298;
  reg [31:0] p5_xor_63300;
  reg [31:0] p5_add_63317;
  reg [31:0] p5_add_63120;
  always_ff @ (posedge clk) begin
    p5_message <= p4_message;
    p5_concat_63072 <= p4_concat_63072;
    p5_add_63143 <= p4_add_63143;
    p5_add_63192 <= p4_add_63192;
    p5_add_63194 <= p4_add_63194;
    p5_add_63273 <= p5_add_63273_comb;
    p5_add_63274 <= p5_add_63274_comb;
    p5_add_63244 <= p4_add_63244;
    p5_add_63297 <= p5_add_63297_comb;
    p5_and_63298 <= p5_and_63298_comb;
    p5_xor_63300 <= p5_xor_63300_comb;
    p5_add_63317 <= p5_add_63317_comb;
    p5_add_63120 <= p4_add_63120;
  end

  // ===== Pipe stage 6:
  wire [31:0] p6_add_63365_comb;
  wire [31:0] p6_add_63368_comb;
  wire [31:0] p6_add_63369_comb;
  wire [31:0] p6_add_63388_comb;
  wire [31:0] p6_add_63370_comb;
  wire [31:0] p6_add_63389_comb;
  wire [31:0] p6_add_63406_comb;
  assign p6_add_63365_comb = {p5_add_63274[5:0] ^ p5_add_63274[10:5] ^ p5_add_63274[24:19], p5_add_63274[31:27] ^ p5_add_63274[4:0] ^ p5_add_63274[18:14], p5_add_63274[26:13] ^ p5_add_63274[31:18] ^ p5_add_63274[13:0], p5_add_63274[12:6] ^ p5_add_63274[17:11] ^ p5_add_63274[31:25]} + (p5_add_63274 & p5_add_63194 ^ ~(p5_add_63274 | ~p5_add_63143));
  assign p6_add_63368_comb = p6_add_63365_comb + 32'h59f1_11f1;
  assign p6_add_63369_comb = p5_concat_63072 + p5_message[351:320];
  assign p6_add_63388_comb = {p5_add_63297[1:0] ^ p5_add_63297[12:11] ^ p5_add_63297[21:20], p5_add_63297[31:21] ^ p5_add_63297[10:0] ^ p5_add_63297[19:9], p5_add_63297[20:12] ^ p5_add_63297[31:23] ^ p5_add_63297[8:0], p5_add_63297[11:2] ^ p5_add_63297[22:13] ^ p5_add_63297[31:22]} + p5_xor_63300;
  assign p6_add_63370_comb = p6_add_63368_comb + p6_add_63369_comb;
  assign p6_add_63389_comb = p5_add_63192 + p6_add_63388_comb;
  assign p6_add_63406_comb = {p5_message[294:292] ^ p5_message[305:303], p5_message[291:288] ^ p5_message[302:299] ^ p5_message[319:316], p5_message[319:309] ^ p5_message[298:288] ^ p5_message[315:305], p5_message[308:295] ^ p5_message[319:306] ^ p5_message[304:291]} + p5_message[351:320];

  // Registers for pipe stage 6:
  reg [511:0] p6_message;
  reg [31:0] p6_add_63143;
  reg [31:0] p6_add_63194;
  reg [31:0] p6_add_63273;
  reg [31:0] p6_add_63274;
  reg [31:0] p6_add_63244;
  reg [31:0] p6_add_63370;
  reg [31:0] p6_add_63297;
  reg [31:0] p6_and_63298;
  reg [31:0] p6_add_63389;
  reg [31:0] p6_add_63406;
  reg [31:0] p6_add_63317;
  reg [31:0] p6_add_63120;
  always_ff @ (posedge clk) begin
    p6_message <= p5_message;
    p6_add_63143 <= p5_add_63143;
    p6_add_63194 <= p5_add_63194;
    p6_add_63273 <= p5_add_63273;
    p6_add_63274 <= p5_add_63274;
    p6_add_63244 <= p5_add_63244;
    p6_add_63370 <= p6_add_63370_comb;
    p6_add_63297 <= p5_add_63297;
    p6_and_63298 <= p5_and_63298;
    p6_add_63389 <= p6_add_63389_comb;
    p6_add_63406 <= p6_add_63406_comb;
    p6_add_63317 <= p5_add_63317;
    p6_add_63120 <= p5_add_63120;
  end

  // ===== Pipe stage 7:
  wire [31:0] p7_add_63433_comb;
  wire [31:0] p7_and_63479_comb;
  wire [29:0] p7_add_63455_comb;
  wire [31:0] p7_add_63483_comb;
  wire [31:0] p7_add_63460_comb;
  wire [31:0] p7_add_63461_comb;
  wire [31:0] p7_add_63484_comb;
  wire [31:0] p7_add_63462_comb;
  assign p7_add_63433_comb = p6_add_63244 + p6_add_63370;
  assign p7_and_63479_comb = p6_add_63389 & p6_add_63297;
  assign p7_add_63455_comb = p6_message[319:290] + 30'h248f_e0a9;
  assign p7_add_63483_comb = {p6_add_63389[1:0] ^ p6_add_63389[12:11] ^ p6_add_63389[21:20], p6_add_63389[31:21] ^ p6_add_63389[10:0] ^ p6_add_63389[19:9], p6_add_63389[20:12] ^ p6_add_63389[31:23] ^ p6_add_63389[8:0], p6_add_63389[11:2] ^ p6_add_63389[22:13] ^ p6_add_63389[31:22]} + (p7_and_63479_comb ^ p6_add_63389 & p6_add_63244 ^ p6_and_63298);
  assign p7_add_63460_comb = {p7_add_63433_comb[5:0] ^ p7_add_63433_comb[10:5] ^ p7_add_63433_comb[24:19], p7_add_63433_comb[31:27] ^ p7_add_63433_comb[4:0] ^ p7_add_63433_comb[18:14], p7_add_63433_comb[26:13] ^ p7_add_63433_comb[31:18] ^ p7_add_63433_comb[13:0], p7_add_63433_comb[12:6] ^ p7_add_63433_comb[17:11] ^ p7_add_63433_comb[31:25]} + p6_add_63143;
  assign p7_add_63461_comb = (p7_add_63433_comb & p6_add_63274 ^ ~(p7_add_63433_comb | ~p6_add_63194)) + {p7_add_63455_comb, p6_message[289:288]};
  assign p7_add_63484_comb = p6_add_63273 + p7_add_63483_comb;
  assign p7_add_63462_comb = p7_add_63460_comb + p7_add_63461_comb;

  // Registers for pipe stage 7:
  reg [511:0] p7_message;
  reg [31:0] p7_add_63194;
  reg [31:0] p7_add_63274;
  reg [31:0] p7_add_63370;
  reg [31:0] p7_add_63433;
  reg [31:0] p7_add_63297;
  reg [31:0] p7_add_63389;
  reg [31:0] p7_and_63479;
  reg [31:0] p7_add_63484;
  reg [31:0] p7_add_63406;
  reg [31:0] p7_add_63317;
  reg [31:0] p7_add_63120;
  reg [31:0] p7_add_63462;
  always_ff @ (posedge clk) begin
    p7_message <= p6_message;
    p7_add_63194 <= p6_add_63194;
    p7_add_63274 <= p6_add_63274;
    p7_add_63370 <= p6_add_63370;
    p7_add_63433 <= p7_add_63433_comb;
    p7_add_63297 <= p6_add_63297;
    p7_add_63389 <= p6_add_63389;
    p7_and_63479 <= p7_and_63479_comb;
    p7_add_63484 <= p7_add_63484_comb;
    p7_add_63406 <= p6_add_63406;
    p7_add_63317 <= p6_add_63317;
    p7_add_63120 <= p6_add_63120;
    p7_add_63462 <= p7_add_63462_comb;
  end

  // ===== Pipe stage 8:
  wire [31:0] p8_add_63511_comb;
  wire [31:0] p8_and_63554_comb;
  wire [31:0] p8_add_63558_comb;
  wire [31:0] p8_add_63533_comb;
  wire [31:0] p8_add_63537_comb;
  wire [31:0] p8_add_63559_comb;
  wire [31:0] p8_add_63536_comb;
  wire [31:0] p8_add_63576_comb;
  assign p8_add_63511_comb = p7_add_63297 + p7_add_63462;
  assign p8_and_63554_comb = p7_add_63484 & p7_add_63389;
  assign p8_add_63558_comb = {p7_add_63484[1:0] ^ p7_add_63484[12:11] ^ p7_add_63484[21:20], p7_add_63484[31:21] ^ p7_add_63484[10:0] ^ p7_add_63484[19:9], p7_add_63484[20:12] ^ p7_add_63484[31:23] ^ p7_add_63484[8:0], p7_add_63484[11:2] ^ p7_add_63484[22:13] ^ p7_add_63484[31:22]} + (p8_and_63554_comb ^ p7_add_63484 & p7_add_63297 ^ p7_and_63479);
  assign p8_add_63533_comb = {p8_add_63511_comb[5:0] ^ p8_add_63511_comb[10:5] ^ p8_add_63511_comb[24:19], p8_add_63511_comb[31:27] ^ p8_add_63511_comb[4:0] ^ p8_add_63511_comb[18:14], p8_add_63511_comb[26:13] ^ p8_add_63511_comb[31:18] ^ p8_add_63511_comb[13:0], p8_add_63511_comb[12:6] ^ p8_add_63511_comb[17:11] ^ p8_add_63511_comb[31:25]} + (p8_add_63511_comb & p7_add_63433 ^ ~(p8_add_63511_comb | ~p7_add_63274));
  assign p8_add_63537_comb = p7_add_63194 + p7_message[287:256];
  assign p8_add_63559_comb = p7_add_63370 + p8_add_63558_comb;
  assign p8_add_63536_comb = p8_add_63533_comb + 32'hab1c_5ed5;
  assign p8_add_63576_comb = {p7_message[230:228] ^ p7_message[241:239], p7_message[227:224] ^ p7_message[238:235] ^ p7_message[255:252], p7_message[255:245] ^ p7_message[234:224] ^ p7_message[251:241], p7_message[244:231] ^ p7_message[255:242] ^ p7_message[240:227]} + p7_message[287:256];

  // Registers for pipe stage 8:
  reg [511:0] p8_message;
  reg [31:0] p8_add_63274;
  reg [31:0] p8_add_63433;
  reg [31:0] p8_add_63511;
  reg [31:0] p8_add_63537;
  reg [31:0] p8_add_63389;
  reg [31:0] p8_add_63484;
  reg [31:0] p8_and_63554;
  reg [31:0] p8_add_63559;
  reg [31:0] p8_add_63536;
  reg [31:0] p8_add_63576;
  reg [31:0] p8_add_63406;
  reg [31:0] p8_add_63317;
  reg [31:0] p8_add_63120;
  reg [31:0] p8_add_63462;
  always_ff @ (posedge clk) begin
    p8_message <= p7_message;
    p8_add_63274 <= p7_add_63274;
    p8_add_63433 <= p7_add_63433;
    p8_add_63511 <= p8_add_63511_comb;
    p8_add_63537 <= p8_add_63537_comb;
    p8_add_63389 <= p7_add_63389;
    p8_add_63484 <= p7_add_63484;
    p8_and_63554 <= p8_and_63554_comb;
    p8_add_63559 <= p8_add_63559_comb;
    p8_add_63536 <= p8_add_63536_comb;
    p8_add_63576 <= p8_add_63576_comb;
    p8_add_63406 <= p7_add_63406;
    p8_add_63317 <= p7_add_63317;
    p8_add_63120 <= p7_add_63120;
    p8_add_63462 <= p7_add_63462;
  end

  // ===== Pipe stage 9:
  wire [31:0] p9_add_63607_comb;
  wire [31:0] p9_add_63608_comb;
  wire [31:0] p9_and_63653_comb;
  wire [28:0] p9_add_63630_comb;
  wire [31:0] p9_add_63657_comb;
  wire [31:0] p9_add_63658_comb;
  wire [31:0] p9_add_63635_comb;
  wire [31:0] p9_add_63636_comb;
  assign p9_add_63607_comb = p8_add_63536 + p8_add_63537;
  assign p9_add_63608_comb = p8_add_63389 + p9_add_63607_comb;
  assign p9_and_63653_comb = p8_add_63559 & p8_add_63484;
  assign p9_add_63630_comb = p8_message[255:227] + 29'h1b00_f553;
  assign p9_add_63657_comb = {p8_add_63559[1:0] ^ p8_add_63559[12:11] ^ p8_add_63559[21:20], p8_add_63559[31:21] ^ p8_add_63559[10:0] ^ p8_add_63559[19:9], p8_add_63559[20:12] ^ p8_add_63559[31:23] ^ p8_add_63559[8:0], p8_add_63559[11:2] ^ p8_add_63559[22:13] ^ p8_add_63559[31:22]} + (p9_and_63653_comb ^ p8_add_63559 & p8_add_63389 ^ p8_and_63554);
  assign p9_add_63658_comb = p8_add_63462 + p9_add_63657_comb;
  assign p9_add_63635_comb = {p9_add_63608_comb[5:0] ^ p9_add_63608_comb[10:5] ^ p9_add_63608_comb[24:19], p9_add_63608_comb[31:27] ^ p9_add_63608_comb[4:0] ^ p9_add_63608_comb[18:14], p9_add_63608_comb[26:13] ^ p9_add_63608_comb[31:18] ^ p9_add_63608_comb[13:0], p9_add_63608_comb[12:6] ^ p9_add_63608_comb[17:11] ^ p9_add_63608_comb[31:25]} + p8_add_63274;
  assign p9_add_63636_comb = (p9_add_63608_comb & p8_add_63511 ^ ~(p9_add_63608_comb | ~p8_add_63433)) + {p9_add_63630_comb, p8_message[226:224]};

  // Registers for pipe stage 9:
  reg [511:0] p9_message;
  reg [31:0] p9_add_63433;
  reg [31:0] p9_add_63511;
  reg [31:0] p9_add_63607;
  reg [31:0] p9_add_63608;
  reg [31:0] p9_add_63484;
  reg [31:0] p9_add_63559;
  reg [31:0] p9_and_63653;
  reg [31:0] p9_add_63658;
  reg [31:0] p9_add_63576;
  reg [31:0] p9_add_63406;
  reg [31:0] p9_add_63317;
  reg [31:0] p9_add_63120;
  reg [31:0] p9_add_63635;
  reg [31:0] p9_add_63636;
  always_ff @ (posedge clk) begin
    p9_message <= p8_message;
    p9_add_63433 <= p8_add_63433;
    p9_add_63511 <= p8_add_63511;
    p9_add_63607 <= p9_add_63607_comb;
    p9_add_63608 <= p9_add_63608_comb;
    p9_add_63484 <= p8_add_63484;
    p9_add_63559 <= p8_add_63559;
    p9_and_63653 <= p9_and_63653_comb;
    p9_add_63658 <= p9_add_63658_comb;
    p9_add_63576 <= p8_add_63576;
    p9_add_63406 <= p8_add_63406;
    p9_add_63317 <= p8_add_63317;
    p9_add_63120 <= p8_add_63120;
    p9_add_63635 <= p9_add_63635_comb;
    p9_add_63636 <= p9_add_63636_comb;
  end

  // ===== Pipe stage 10:
  wire [31:0] p10_add_63689_comb;
  wire [31:0] p10_add_63690_comb;
  wire [31:0] p10_and_63729_comb;
  wire [31:0] p10_add_63733_comb;
  wire [31:0] p10_add_63712_comb;
  wire [31:0] p10_add_63734_comb;
  assign p10_add_63689_comb = p9_add_63635 + p9_add_63636;
  assign p10_add_63690_comb = p9_add_63484 + p10_add_63689_comb;
  assign p10_and_63729_comb = p9_add_63658 & p9_add_63559;
  assign p10_add_63733_comb = {p9_add_63658[1:0] ^ p9_add_63658[12:11] ^ p9_add_63658[21:20], p9_add_63658[31:21] ^ p9_add_63658[10:0] ^ p9_add_63658[19:9], p9_add_63658[20:12] ^ p9_add_63658[31:23] ^ p9_add_63658[8:0], p9_add_63658[11:2] ^ p9_add_63658[22:13] ^ p9_add_63658[31:22]} + (p10_and_63729_comb ^ p9_add_63658 & p9_add_63484 ^ p9_and_63653);
  assign p10_add_63712_comb = {p10_add_63690_comb[5:0] ^ p10_add_63690_comb[10:5] ^ p10_add_63690_comb[24:19], p10_add_63690_comb[31:27] ^ p10_add_63690_comb[4:0] ^ p10_add_63690_comb[18:14], p10_add_63690_comb[26:13] ^ p10_add_63690_comb[31:18] ^ p10_add_63690_comb[13:0], p10_add_63690_comb[12:6] ^ p10_add_63690_comb[17:11] ^ p10_add_63690_comb[31:25]} + (p10_add_63690_comb & p9_add_63608 ^ ~(p10_add_63690_comb | ~p9_add_63511));
  assign p10_add_63734_comb = p9_add_63607 + p10_add_63733_comb;

  // Registers for pipe stage 10:
  reg [511:0] p10_message;
  reg [31:0] p10_add_63433;
  reg [31:0] p10_add_63511;
  reg [31:0] p10_add_63608;
  reg [31:0] p10_add_63690;
  reg [31:0] p10_add_63712;
  reg [31:0] p10_add_63559;
  reg [31:0] p10_add_63658;
  reg [31:0] p10_and_63729;
  reg [31:0] p10_add_63734;
  reg [31:0] p10_add_63576;
  reg [31:0] p10_add_63406;
  reg [31:0] p10_add_63317;
  reg [31:0] p10_add_63120;
  reg [31:0] p10_add_63689;
  always_ff @ (posedge clk) begin
    p10_message <= p9_message;
    p10_add_63433 <= p9_add_63433;
    p10_add_63511 <= p9_add_63511;
    p10_add_63608 <= p9_add_63608;
    p10_add_63690 <= p10_add_63690_comb;
    p10_add_63712 <= p10_add_63712_comb;
    p10_add_63559 <= p9_add_63559;
    p10_add_63658 <= p9_add_63658;
    p10_and_63729 <= p10_and_63729_comb;
    p10_add_63734 <= p10_add_63734_comb;
    p10_add_63576 <= p9_add_63576;
    p10_add_63406 <= p9_add_63406;
    p10_add_63317 <= p9_add_63317;
    p10_add_63120 <= p9_add_63120;
    p10_add_63689 <= p10_add_63689_comb;
  end

  // ===== Pipe stage 11:
  wire [31:0] p11_and_63790_comb;
  wire [31:0] p11_add_63767_comb;
  wire [31:0] p11_add_63768_comb;
  wire [31:0] p11_add_63769_comb;
  wire [31:0] p11_add_63794_comb;
  wire [31:0] p11_add_63829_comb;
  wire [31:0] p11_add_63830_comb;
  wire [31:0] p11_add_63770_comb;
  wire [30:0] p11_add_63773_comb;
  wire [31:0] p11_add_63795_comb;
  wire [31:0] p11_add_63848_comb;
  wire [31:0] p11_add_63831_comb;
  assign p11_and_63790_comb = p10_add_63734 & p10_add_63658;
  assign p11_add_63767_comb = p10_add_63712 + 32'h1283_5b01;
  assign p11_add_63768_comb = p10_add_63433 + p10_message[223:192];
  assign p11_add_63769_comb = p11_add_63767_comb + p11_add_63768_comb;
  assign p11_add_63794_comb = {p10_add_63734[1:0] ^ p10_add_63734[12:11] ^ p10_add_63734[21:20], p10_add_63734[31:21] ^ p10_add_63734[10:0] ^ p10_add_63734[19:9], p10_add_63734[20:12] ^ p10_add_63734[31:23] ^ p10_add_63734[8:0], p10_add_63734[11:2] ^ p10_add_63734[22:13] ^ p10_add_63734[31:22]} + (p11_and_63790_comb ^ p10_add_63734 & p10_add_63559 ^ p10_and_63729);
  assign p11_add_63829_comb = {p10_message[454:452] ^ p10_message[465:463], p10_message[451:448] ^ p10_message[462:459] ^ p10_message[479:476], p10_message[479:469] ^ p10_message[458:448] ^ p10_message[475:465], p10_message[468:455] ^ p10_message[479:466] ^ p10_message[464:451]} + p10_message[511:480];
  assign p11_add_63830_comb = p10_message[223:192] + {p10_message[48:39] ^ p10_message[50:41], p10_message[38:32] ^ p10_message[40:34] ^ p10_message[63:57], p10_message[63:62] ^ p10_message[33:32] ^ p10_message[56:55], p10_message[61:49] ^ p10_message[63:51] ^ p10_message[54:42]};
  assign p11_add_63770_comb = p10_add_63559 + p11_add_63769_comb;
  assign p11_add_63773_comb = p10_message[191:161] + 31'h1218_c2df;
  assign p11_add_63795_comb = p10_add_63689 + p11_add_63794_comb;
  assign p11_add_63848_comb = {p10_message[166:164] ^ p10_message[177:175], p10_message[163:160] ^ p10_message[174:171] ^ p10_message[191:188], p10_message[191:181] ^ p10_message[170:160] ^ p10_message[187:177], p10_message[180:167] ^ p10_message[191:178] ^ p10_message[176:163]} + p10_message[223:192];
  assign p11_add_63831_comb = p11_add_63829_comb + p11_add_63830_comb;

  // Registers for pipe stage 11:
  reg [511:0] p11_message;
  reg [31:0] p11_add_63511;
  reg [31:0] p11_add_63608;
  reg [31:0] p11_add_63690;
  reg [31:0] p11_add_63769;
  reg [31:0] p11_add_63770;
  reg [30:0] p11_add_63773;
  reg [31:0] p11_add_63658;
  reg [31:0] p11_add_63734;
  reg [31:0] p11_and_63790;
  reg [31:0] p11_add_63795;
  reg [31:0] p11_add_63848;
  reg [31:0] p11_add_63576;
  reg [31:0] p11_add_63406;
  reg [31:0] p11_add_63317;
  reg [31:0] p11_add_63120;
  reg [31:0] p11_add_63831;
  always_ff @ (posedge clk) begin
    p11_message <= p10_message;
    p11_add_63511 <= p10_add_63511;
    p11_add_63608 <= p10_add_63608;
    p11_add_63690 <= p10_add_63690;
    p11_add_63769 <= p11_add_63769_comb;
    p11_add_63770 <= p11_add_63770_comb;
    p11_add_63773 <= p11_add_63773_comb;
    p11_add_63658 <= p10_add_63658;
    p11_add_63734 <= p10_add_63734;
    p11_and_63790 <= p11_and_63790_comb;
    p11_add_63795 <= p11_add_63795_comb;
    p11_add_63848 <= p11_add_63848_comb;
    p11_add_63576 <= p10_add_63576;
    p11_add_63406 <= p10_add_63406;
    p11_add_63317 <= p10_add_63317;
    p11_add_63120 <= p10_add_63120;
    p11_add_63831 <= p11_add_63831_comb;
  end

  // ===== Pipe stage 12:
  wire [31:0] p12_add_64002_comb;
  wire [31:0] p12_add_63983_comb;
  wire [31:0] p12_add_63984_comb;
  wire [31:0] p12_add_64003_comb;
  wire [31:0] p12_add_63985_comb;
  wire [31:0] p12_and_63935_comb;
  wire [31:0] p12_add_63906_comb;
  wire [31:0] p12_add_63907_comb;
  wire [31:0] p12_add_63908_comb;
  wire [29:0] p12_add_63914_comb;
  wire [30:0] p12_add_63937_comb;
  wire [31:0] p12_add_63942_comb;
  wire [29:0] p12_add_63947_comb;
  wire [31:0] p12_bit_slice_63944_comb;
  wire [31:0] p12_add_63909_comb;
  wire [31:0] p12_add_63911_comb;
  wire [31:0] p12_concat_63916_comb;
  wire [31:0] p12_concat_63941_comb;
  wire [31:0] p12_add_63943_comb;
  wire [31:0] p12_concat_63949_comb;
  wire [31:0] p12_bit_slice_64075_comb;
  wire [31:0] p12_add_64179_comb;
  wire [31:0] p12_add_64162_comb;
  wire [31:0] p12_add_64145_comb;
  wire [31:0] p12_add_64128_comb;
  wire [31:0] p12_add_64111_comb;
  wire [31:0] p12_add_64094_comb;
  wire [31:0] p12_add_64076_comb;
  wire [31:0] p12_add_64057_comb;
  wire [31:0] p12_add_64038_comb;
  wire [31:0] p12_add_64039_comb;
  assign p12_add_64002_comb = p11_message[159:128] + {p11_add_63831[16:7] ^ p11_add_63831[18:9], p11_add_63831[6:0] ^ p11_add_63831[8:2] ^ p11_add_63831[31:25], p11_add_63831[31:30] ^ p11_add_63831[1:0] ^ p11_add_63831[24:23], p11_add_63831[29:17] ^ p11_add_63831[31:19] ^ p11_add_63831[22:10]};
  assign p12_add_63983_comb = {p11_message[422:420] ^ p11_message[433:431], p11_message[419:416] ^ p11_message[430:427] ^ p11_message[447:444], p11_message[447:437] ^ p11_message[426:416] ^ p11_message[443:433], p11_message[436:423] ^ p11_message[447:434] ^ p11_message[432:419]} + p11_message[479:448];
  assign p12_add_63984_comb = p11_message[191:160] + {p11_message[16:7] ^ p11_message[18:9], p11_message[6:0] ^ p11_message[8:2] ^ p11_message[31:25], p11_message[31:30] ^ p11_message[1:0] ^ p11_message[24:23], p11_message[29:17] ^ p11_message[31:19] ^ p11_message[22:10]};
  assign p12_add_64003_comb = p11_add_63120 + p12_add_64002_comb;
  assign p12_add_63985_comb = p12_add_63983_comb + p12_add_63984_comb;
  assign p12_and_63935_comb = p11_add_63795 & p11_add_63734;
  assign p12_add_63906_comb = {p11_add_63770[5:0] ^ p11_add_63770[10:5] ^ p11_add_63770[24:19], p11_add_63770[31:27] ^ p11_add_63770[4:0] ^ p11_add_63770[18:14], p11_add_63770[26:13] ^ p11_add_63770[31:18] ^ p11_add_63770[13:0], p11_add_63770[12:6] ^ p11_add_63770[17:11] ^ p11_add_63770[31:25]} + p11_add_63511;
  assign p12_add_63907_comb = (p11_add_63770 & p11_add_63690 ^ ~(p11_add_63770 | ~p11_add_63608)) + {p11_add_63773, p11_message[160]};
  assign p12_add_63908_comb = p12_add_63906_comb + p12_add_63907_comb;
  assign p12_add_63914_comb = p11_message[127:98] + 30'h1caf_975d;
  assign p12_add_63937_comb = p11_message[95:65] + 31'h406f_58ff;
  assign p12_add_63942_comb = {p11_add_63795[1:0] ^ p11_add_63795[12:11] ^ p11_add_63795[21:20], p11_add_63795[31:21] ^ p11_add_63795[10:0] ^ p11_add_63795[19:9], p11_add_63795[20:12] ^ p11_add_63795[31:23] ^ p11_add_63795[8:0], p11_add_63795[11:2] ^ p11_add_63795[22:13] ^ p11_add_63795[31:22]} + (p12_and_63935_comb ^ p11_add_63795 & p11_add_63658 ^ p11_and_63790);
  assign p12_add_63947_comb = p11_message[31:2] + 30'h3066_fc5d;
  assign p12_bit_slice_63944_comb = p11_message[63:32];
  assign p12_add_63909_comb = p11_add_63658 + p12_add_63908_comb;
  assign p12_add_63911_comb = p11_add_63608 + p11_message[159:128];
  assign p12_concat_63916_comb = {p12_add_63914_comb, p11_message[97:96]};
  assign p12_concat_63941_comb = {p12_add_63937_comb, p11_message[64]};
  assign p12_add_63943_comb = p11_add_63769 + p12_add_63942_comb;
  assign p12_concat_63949_comb = {p12_add_63947_comb, p11_message[1:0]};
  assign p12_bit_slice_64075_comb = p11_message[31:0];
  assign p12_add_64179_comb = {p11_message[6:4] ^ p11_message[17:15], p11_message[3:0] ^ p11_message[14:11] ^ p11_message[31:28], p11_message[31:21] ^ p11_message[10:0] ^ p11_message[27:17], p11_message[20:7] ^ p11_message[31:18] ^ p11_message[16:3]} + p12_bit_slice_63944_comb;
  assign p12_add_64162_comb = {p11_message[38:36] ^ p11_message[49:47], p11_message[35:32] ^ p11_message[46:43] ^ p11_message[63:60], p11_message[63:53] ^ p11_message[42:32] ^ p11_message[59:49], p11_message[52:39] ^ p11_message[63:50] ^ p11_message[48:35]} + p11_message[95:64];
  assign p12_add_64145_comb = {p11_message[70:68] ^ p11_message[81:79], p11_message[67:64] ^ p11_message[78:75] ^ p11_message[95:92], p11_message[95:85] ^ p11_message[74:64] ^ p11_message[91:81], p11_message[84:71] ^ p11_message[95:82] ^ p11_message[80:67]} + p11_message[127:96];
  assign p12_add_64128_comb = {p11_message[102:100] ^ p11_message[113:111], p11_message[99:96] ^ p11_message[110:107] ^ p11_message[127:124], p11_message[127:117] ^ p11_message[106:96] ^ p11_message[123:113], p11_message[116:103] ^ p11_message[127:114] ^ p11_message[112:99]} + p11_message[159:128];
  assign p12_add_64111_comb = {p11_message[134:132] ^ p11_message[145:143], p11_message[131:128] ^ p11_message[142:139] ^ p11_message[159:156], p11_message[159:149] ^ p11_message[138:128] ^ p11_message[155:145], p11_message[148:135] ^ p11_message[159:146] ^ p11_message[144:131]} + p11_message[191:160];
  assign p12_add_64094_comb = {p11_message[198:196] ^ p11_message[209:207], p11_message[195:192] ^ p11_message[206:203] ^ p11_message[223:220], p11_message[223:213] ^ p11_message[202:192] ^ p11_message[219:209], p11_message[212:199] ^ p11_message[223:210] ^ p11_message[208:195]} + p11_message[255:224];
  assign p12_add_64076_comb = {p11_message[262:260] ^ p11_message[273:271], p11_message[259:256] ^ p11_message[270:267] ^ p11_message[287:284], p11_message[287:277] ^ p11_message[266:256] ^ p11_message[283:273], p11_message[276:263] ^ p11_message[287:274] ^ p11_message[272:259]} + p11_message[319:288];
  assign p12_add_64057_comb = p11_message[95:64] + {p12_add_64003_comb[16:7] ^ p12_add_64003_comb[18:9], p12_add_64003_comb[6:0] ^ p12_add_64003_comb[8:2] ^ p12_add_64003_comb[31:25], p12_add_64003_comb[31:30] ^ p12_add_64003_comb[1:0] ^ p12_add_64003_comb[24:23], p12_add_64003_comb[29:17] ^ p12_add_64003_comb[31:19] ^ p12_add_64003_comb[22:10]};
  assign p12_add_64038_comb = {p11_message[358:356] ^ p11_message[369:367], p11_message[355:352] ^ p11_message[366:363] ^ p11_message[383:380], p11_message[383:373] ^ p11_message[362:352] ^ p11_message[379:369], p11_message[372:359] ^ p11_message[383:370] ^ p11_message[368:355]} + p11_message[415:384];
  assign p12_add_64039_comb = p11_message[127:96] + {p12_add_63985_comb[16:7] ^ p12_add_63985_comb[18:9], p12_add_63985_comb[6:0] ^ p12_add_63985_comb[8:2] ^ p12_add_63985_comb[31:25], p12_add_63985_comb[31:30] ^ p12_add_63985_comb[1:0] ^ p12_add_63985_comb[24:23], p12_add_63985_comb[29:17] ^ p12_add_63985_comb[31:19] ^ p12_add_63985_comb[22:10]};

  // Registers for pipe stage 12:
  reg [31:0] p12_add_63690;
  reg [31:0] p12_add_63770;
  reg [31:0] p12_add_63909;
  reg [31:0] p12_add_63911;
  reg [31:0] p12_add_63734;
  reg [31:0] p12_concat_63916;
  reg [31:0] p12_add_63795;
  reg [31:0] p12_and_63935;
  reg [31:0] p12_concat_63941;
  reg [31:0] p12_add_63943;
  reg [31:0] p12_bit_slice_63944;
  reg [31:0] p12_concat_63949;
  reg [31:0] p12_bit_slice_64075;
  reg [31:0] p12_add_64179;
  reg [31:0] p12_add_64162;
  reg [31:0] p12_add_64145;
  reg [31:0] p12_add_64128;
  reg [31:0] p12_add_64111;
  reg [31:0] p12_add_63848;
  reg [31:0] p12_add_64094;
  reg [31:0] p12_add_63576;
  reg [31:0] p12_add_64076;
  reg [31:0] p12_add_63406;
  reg [31:0] p12_add_63317;
  reg [31:0] p12_add_64057;
  reg [31:0] p12_add_64038;
  reg [31:0] p12_add_64039;
  reg [31:0] p12_add_64003;
  reg [31:0] p12_add_63985;
  reg [31:0] p12_add_63831;
  reg [31:0] p12_add_63908;
  always_ff @ (posedge clk) begin
    p12_add_63690 <= p11_add_63690;
    p12_add_63770 <= p11_add_63770;
    p12_add_63909 <= p12_add_63909_comb;
    p12_add_63911 <= p12_add_63911_comb;
    p12_add_63734 <= p11_add_63734;
    p12_concat_63916 <= p12_concat_63916_comb;
    p12_add_63795 <= p11_add_63795;
    p12_and_63935 <= p12_and_63935_comb;
    p12_concat_63941 <= p12_concat_63941_comb;
    p12_add_63943 <= p12_add_63943_comb;
    p12_bit_slice_63944 <= p12_bit_slice_63944_comb;
    p12_concat_63949 <= p12_concat_63949_comb;
    p12_bit_slice_64075 <= p12_bit_slice_64075_comb;
    p12_add_64179 <= p12_add_64179_comb;
    p12_add_64162 <= p12_add_64162_comb;
    p12_add_64145 <= p12_add_64145_comb;
    p12_add_64128 <= p12_add_64128_comb;
    p12_add_64111 <= p12_add_64111_comb;
    p12_add_63848 <= p11_add_63848;
    p12_add_64094 <= p12_add_64094_comb;
    p12_add_63576 <= p11_add_63576;
    p12_add_64076 <= p12_add_64076_comb;
    p12_add_63406 <= p11_add_63406;
    p12_add_63317 <= p11_add_63317;
    p12_add_64057 <= p12_add_64057_comb;
    p12_add_64038 <= p12_add_64038_comb;
    p12_add_64039 <= p12_add_64039_comb;
    p12_add_64003 <= p12_add_64003_comb;
    p12_add_63985 <= p12_add_63985_comb;
    p12_add_63831 <= p11_add_63831;
    p12_add_63908 <= p12_add_63908_comb;
  end

  // ===== Pipe stage 13:
  wire [31:0] p13_add_64290_comb;
  wire [31:0] p13_and_64283_comb;
  wire [31:0] p13_add_64263_comb;
  wire [31:0] p13_add_64265_comb;
  wire [31:0] p13_add_64287_comb;
  wire [31:0] p13_add_64307_comb;
  wire [31:0] p13_add_64266_comb;
  wire [31:0] p13_add_64288_comb;
  wire [31:0] p13_add_64325_comb;
  wire [31:0] p13_add_64308_comb;
  wire [31:0] p13_add_64289_comb;
  assign p13_add_64290_comb = p12_add_63317 + p12_add_64057;
  assign p13_and_64283_comb = p12_add_63943 & p12_add_63795;
  assign p13_add_64263_comb = {p12_add_63909[5:0] ^ p12_add_63909[10:5] ^ p12_add_63909[24:19], p12_add_63909[31:27] ^ p12_add_63909[4:0] ^ p12_add_63909[18:14], p12_add_63909[26:13] ^ p12_add_63909[31:18] ^ p12_add_63909[13:0], p12_add_63909[12:6] ^ p12_add_63909[17:11] ^ p12_add_63909[31:25]} + (p12_add_63909 & p12_add_63770 ^ ~(p12_add_63909 | ~p12_add_63690));
  assign p13_add_64265_comb = p13_add_64263_comb + 32'h550c_7dc3;
  assign p13_add_64287_comb = {p12_add_63943[1:0] ^ p12_add_63943[12:11] ^ p12_add_63943[21:20], p12_add_63943[31:21] ^ p12_add_63943[10:0] ^ p12_add_63943[19:9], p12_add_63943[20:12] ^ p12_add_63943[31:23] ^ p12_add_63943[8:0], p12_add_63943[11:2] ^ p12_add_63943[22:13] ^ p12_add_63943[31:22]} + (p13_and_64283_comb ^ p12_add_63943 & p12_add_63734 ^ p12_and_63935);
  assign p13_add_64307_comb = p12_bit_slice_64075 + {p13_add_64290_comb[16:7] ^ p13_add_64290_comb[18:9], p13_add_64290_comb[6:0] ^ p13_add_64290_comb[8:2] ^ p13_add_64290_comb[31:25], p13_add_64290_comb[31:30] ^ p13_add_64290_comb[1:0] ^ p13_add_64290_comb[24:23], p13_add_64290_comb[29:17] ^ p13_add_64290_comb[31:19] ^ p13_add_64290_comb[22:10]};
  assign p13_add_64266_comb = p13_add_64265_comb + p12_add_63911;
  assign p13_add_64288_comb = p12_add_63908 + p13_add_64287_comb;
  assign p13_add_64325_comb = {p12_add_63831[6:4] ^ p12_add_63831[17:15], p12_add_63831[3:0] ^ p12_add_63831[14:11] ^ p12_add_63831[31:28], p12_add_63831[31:21] ^ p12_add_63831[10:0] ^ p12_add_63831[27:17], p12_add_63831[20:7] ^ p12_add_63831[31:18] ^ p12_add_63831[16:3]} + p12_bit_slice_64075;
  assign p13_add_64308_comb = p12_add_64076 + p13_add_64307_comb;
  assign p13_add_64289_comb = p12_add_64038 + p12_add_64039;

  // Registers for pipe stage 13:
  reg [31:0] p13_add_63690;
  reg [31:0] p13_add_63770;
  reg [31:0] p13_add_63909;
  reg [31:0] p13_add_63734;
  reg [31:0] p13_add_64266;
  reg [31:0] p13_concat_63916;
  reg [31:0] p13_add_63795;
  reg [31:0] p13_concat_63941;
  reg [31:0] p13_add_63943;
  reg [31:0] p13_and_64283;
  reg [31:0] p13_bit_slice_63944;
  reg [31:0] p13_add_64288;
  reg [31:0] p13_concat_63949;
  reg [31:0] p13_add_64325;
  reg [31:0] p13_add_64179;
  reg [31:0] p13_add_64162;
  reg [31:0] p13_add_64145;
  reg [31:0] p13_add_64128;
  reg [31:0] p13_add_64111;
  reg [31:0] p13_add_63848;
  reg [31:0] p13_add_64094;
  reg [31:0] p13_add_63576;
  reg [31:0] p13_add_64308;
  reg [31:0] p13_add_63406;
  reg [31:0] p13_add_64290;
  reg [31:0] p13_add_64289;
  reg [31:0] p13_add_64003;
  reg [31:0] p13_add_63985;
  reg [31:0] p13_add_63831;
  always_ff @ (posedge clk) begin
    p13_add_63690 <= p12_add_63690;
    p13_add_63770 <= p12_add_63770;
    p13_add_63909 <= p12_add_63909;
    p13_add_63734 <= p12_add_63734;
    p13_add_64266 <= p13_add_64266_comb;
    p13_concat_63916 <= p12_concat_63916;
    p13_add_63795 <= p12_add_63795;
    p13_concat_63941 <= p12_concat_63941;
    p13_add_63943 <= p12_add_63943;
    p13_and_64283 <= p13_and_64283_comb;
    p13_bit_slice_63944 <= p12_bit_slice_63944;
    p13_add_64288 <= p13_add_64288_comb;
    p13_concat_63949 <= p12_concat_63949;
    p13_add_64325 <= p13_add_64325_comb;
    p13_add_64179 <= p12_add_64179;
    p13_add_64162 <= p12_add_64162;
    p13_add_64145 <= p12_add_64145;
    p13_add_64128 <= p12_add_64128;
    p13_add_64111 <= p12_add_64111;
    p13_add_63848 <= p12_add_63848;
    p13_add_64094 <= p12_add_64094;
    p13_add_63576 <= p12_add_63576;
    p13_add_64308 <= p13_add_64308_comb;
    p13_add_63406 <= p12_add_63406;
    p13_add_64290 <= p13_add_64290_comb;
    p13_add_64289 <= p13_add_64289_comb;
    p13_add_64003 <= p12_add_64003;
    p13_add_63985 <= p12_add_63985;
    p13_add_63831 <= p12_add_63831;
  end

  // ===== Pipe stage 14:
  wire [31:0] p14_add_64384_comb;
  wire [31:0] p14_and_64425_comb;
  wire [31:0] p14_add_64429_comb;
  wire [31:0] p14_add_64406_comb;
  wire [31:0] p14_add_64407_comb;
  wire [31:0] p14_add_64430_comb;
  wire [31:0] p14_add_64408_comb;
  assign p14_add_64384_comb = p13_add_63734 + p13_add_64266;
  assign p14_and_64425_comb = p13_add_64288 & p13_add_63943;
  assign p14_add_64429_comb = {p13_add_64288[1:0] ^ p13_add_64288[12:11] ^ p13_add_64288[21:20], p13_add_64288[31:21] ^ p13_add_64288[10:0] ^ p13_add_64288[19:9], p13_add_64288[20:12] ^ p13_add_64288[31:23] ^ p13_add_64288[8:0], p13_add_64288[11:2] ^ p13_add_64288[22:13] ^ p13_add_64288[31:22]} + (p14_and_64425_comb ^ p13_add_64288 & p13_add_63795 ^ p13_and_64283);
  assign p14_add_64406_comb = {p14_add_64384_comb[5:0] ^ p14_add_64384_comb[10:5] ^ p14_add_64384_comb[24:19], p14_add_64384_comb[31:27] ^ p14_add_64384_comb[4:0] ^ p14_add_64384_comb[18:14], p14_add_64384_comb[26:13] ^ p14_add_64384_comb[31:18] ^ p14_add_64384_comb[13:0], p14_add_64384_comb[12:6] ^ p14_add_64384_comb[17:11] ^ p14_add_64384_comb[31:25]} + p13_add_63690;
  assign p14_add_64407_comb = (p14_add_64384_comb & p13_add_63909 ^ ~(p14_add_64384_comb | ~p13_add_63770)) + p13_concat_63916;
  assign p14_add_64430_comb = p13_add_64266 + p14_add_64429_comb;
  assign p14_add_64408_comb = p14_add_64406_comb + p14_add_64407_comb;

  // Registers for pipe stage 14:
  reg [31:0] p14_add_63770;
  reg [31:0] p14_add_63909;
  reg [31:0] p14_add_64384;
  reg [31:0] p14_add_63795;
  reg [31:0] p14_concat_63941;
  reg [31:0] p14_add_63943;
  reg [31:0] p14_bit_slice_63944;
  reg [31:0] p14_add_64288;
  reg [31:0] p14_and_64425;
  reg [31:0] p14_concat_63949;
  reg [31:0] p14_add_64430;
  reg [31:0] p14_add_64325;
  reg [31:0] p14_add_64179;
  reg [31:0] p14_add_64162;
  reg [31:0] p14_add_64145;
  reg [31:0] p14_add_64128;
  reg [31:0] p14_add_64111;
  reg [31:0] p14_add_63848;
  reg [31:0] p14_add_64094;
  reg [31:0] p14_add_63576;
  reg [31:0] p14_add_64308;
  reg [31:0] p14_add_63406;
  reg [31:0] p14_add_64290;
  reg [31:0] p14_add_64289;
  reg [31:0] p14_add_64003;
  reg [31:0] p14_add_63985;
  reg [31:0] p14_add_63831;
  reg [31:0] p14_add_64408;
  always_ff @ (posedge clk) begin
    p14_add_63770 <= p13_add_63770;
    p14_add_63909 <= p13_add_63909;
    p14_add_64384 <= p14_add_64384_comb;
    p14_add_63795 <= p13_add_63795;
    p14_concat_63941 <= p13_concat_63941;
    p14_add_63943 <= p13_add_63943;
    p14_bit_slice_63944 <= p13_bit_slice_63944;
    p14_add_64288 <= p13_add_64288;
    p14_and_64425 <= p14_and_64425_comb;
    p14_concat_63949 <= p13_concat_63949;
    p14_add_64430 <= p14_add_64430_comb;
    p14_add_64325 <= p13_add_64325;
    p14_add_64179 <= p13_add_64179;
    p14_add_64162 <= p13_add_64162;
    p14_add_64145 <= p13_add_64145;
    p14_add_64128 <= p13_add_64128;
    p14_add_64111 <= p13_add_64111;
    p14_add_63848 <= p13_add_63848;
    p14_add_64094 <= p13_add_64094;
    p14_add_63576 <= p13_add_63576;
    p14_add_64308 <= p13_add_64308;
    p14_add_63406 <= p13_add_63406;
    p14_add_64290 <= p13_add_64290;
    p14_add_64289 <= p13_add_64289;
    p14_add_64003 <= p13_add_64003;
    p14_add_63985 <= p13_add_63985;
    p14_add_63831 <= p13_add_63831;
    p14_add_64408 <= p14_add_64408_comb;
  end

  // ===== Pipe stage 15:
  wire [31:0] p15_add_64487_comb;
  wire [1:0] p15_bit_slice_64535_comb;
  wire [31:0] p15_and_64529_comb;
  wire [31:0] p15_add_64533_comb;
  wire [31:0] p15_add_64551_comb;
  wire [31:0] p15_add_64509_comb;
  wire [31:0] p15_add_64510_comb;
  wire [31:0] p15_add_64512_comb;
  wire [31:0] p15_add_64534_comb;
  wire [31:0] p15_add_64552_comb;
  wire [31:0] p15_add_64511_comb;
  assign p15_add_64487_comb = p14_add_63795 + p14_add_64408;
  assign p15_bit_slice_64535_comb = p14_add_64289[1:0];
  assign p15_and_64529_comb = p14_add_64430 & p14_add_64288;
  assign p15_add_64533_comb = {p14_add_64430[1:0] ^ p14_add_64430[12:11] ^ p14_add_64430[21:20], p14_add_64430[31:21] ^ p14_add_64430[10:0] ^ p14_add_64430[19:9], p14_add_64430[20:12] ^ p14_add_64430[31:23] ^ p14_add_64430[8:0], p14_add_64430[11:2] ^ p14_add_64430[22:13] ^ p14_add_64430[31:22]} + (p15_and_64529_comb ^ p14_add_64430 & p14_add_63943 ^ p14_and_64425);
  assign p15_add_64551_comb = p14_bit_slice_63944 + {p14_add_64289[16:7] ^ p14_add_64289[18:9], p14_add_64289[6:0] ^ p14_add_64289[8:2] ^ p14_add_64289[31:25], p14_add_64289[31:30] ^ p15_bit_slice_64535_comb ^ p14_add_64289[24:23], p14_add_64289[29:17] ^ p14_add_64289[31:19] ^ p14_add_64289[22:10]};
  assign p15_add_64509_comb = {p15_add_64487_comb[5:0] ^ p15_add_64487_comb[10:5] ^ p15_add_64487_comb[24:19], p15_add_64487_comb[31:27] ^ p15_add_64487_comb[4:0] ^ p15_add_64487_comb[18:14], p15_add_64487_comb[26:13] ^ p15_add_64487_comb[31:18] ^ p15_add_64487_comb[13:0], p15_add_64487_comb[12:6] ^ p15_add_64487_comb[17:11] ^ p15_add_64487_comb[31:25]} + p14_add_63770;
  assign p15_add_64510_comb = (p15_add_64487_comb & p14_add_64384 ^ ~(p15_add_64487_comb | ~p14_add_63909)) + p14_concat_63941;
  assign p15_add_64512_comb = p14_add_63909 + p14_bit_slice_63944;
  assign p15_add_64534_comb = p14_add_64408 + p15_add_64533_comb;
  assign p15_add_64552_comb = p14_add_63406 + p15_add_64551_comb;
  assign p15_add_64511_comb = p15_add_64509_comb + p15_add_64510_comb;

  // Registers for pipe stage 15:
  reg [31:0] p15_add_64384;
  reg [31:0] p15_add_64487;
  reg [31:0] p15_add_63943;
  reg [31:0] p15_add_64512;
  reg [31:0] p15_add_64288;
  reg [31:0] p15_concat_63949;
  reg [31:0] p15_add_64430;
  reg [31:0] p15_and_64529;
  reg [31:0] p15_add_64534;
  reg [1:0] p15_bit_slice_64535;
  reg [31:0] p15_add_64325;
  reg [31:0] p15_add_64179;
  reg [31:0] p15_add_64162;
  reg [31:0] p15_add_64145;
  reg [31:0] p15_add_64128;
  reg [31:0] p15_add_64111;
  reg [31:0] p15_add_63848;
  reg [31:0] p15_add_64094;
  reg [31:0] p15_add_63576;
  reg [31:0] p15_add_64308;
  reg [31:0] p15_add_64552;
  reg [31:0] p15_add_64290;
  reg [31:0] p15_add_64289;
  reg [31:0] p15_add_64003;
  reg [31:0] p15_add_63985;
  reg [31:0] p15_add_63831;
  reg [31:0] p15_add_64511;
  always_ff @ (posedge clk) begin
    p15_add_64384 <= p14_add_64384;
    p15_add_64487 <= p15_add_64487_comb;
    p15_add_63943 <= p14_add_63943;
    p15_add_64512 <= p15_add_64512_comb;
    p15_add_64288 <= p14_add_64288;
    p15_concat_63949 <= p14_concat_63949;
    p15_add_64430 <= p14_add_64430;
    p15_and_64529 <= p15_and_64529_comb;
    p15_add_64534 <= p15_add_64534_comb;
    p15_bit_slice_64535 <= p15_bit_slice_64535_comb;
    p15_add_64325 <= p14_add_64325;
    p15_add_64179 <= p14_add_64179;
    p15_add_64162 <= p14_add_64162;
    p15_add_64145 <= p14_add_64145;
    p15_add_64128 <= p14_add_64128;
    p15_add_64111 <= p14_add_64111;
    p15_add_63848 <= p14_add_63848;
    p15_add_64094 <= p14_add_64094;
    p15_add_63576 <= p14_add_63576;
    p15_add_64308 <= p14_add_64308;
    p15_add_64552 <= p15_add_64552_comb;
    p15_add_64290 <= p14_add_64290;
    p15_add_64289 <= p14_add_64289;
    p15_add_64003 <= p14_add_64003;
    p15_add_63985 <= p14_add_63985;
    p15_add_63831 <= p14_add_63831;
    p15_add_64511 <= p15_add_64511_comb;
  end

  // ===== Pipe stage 16:
  wire [31:0] p16_add_64607_comb;
  wire [31:0] p16_and_64648_comb;
  wire [31:0] p16_add_64652_comb;
  wire [31:0] p16_add_64629_comb;
  wire [31:0] p16_add_64670_comb;
  wire [31:0] p16_add_64653_comb;
  wire [31:0] p16_add_64631_comb;
  wire [31:0] p16_add_64671_comb;
  assign p16_add_64607_comb = p15_add_63943 + p15_add_64511;
  assign p16_and_64648_comb = p15_add_64534 & p15_add_64430;
  assign p16_add_64652_comb = {p15_add_64534[1:0] ^ p15_add_64534[12:11] ^ p15_add_64534[21:20], p15_add_64534[31:21] ^ p15_add_64534[10:0] ^ p15_add_64534[19:9], p15_add_64534[20:12] ^ p15_add_64534[31:23] ^ p15_add_64534[8:0], p15_add_64534[11:2] ^ p15_add_64534[22:13] ^ p15_add_64534[31:22]} + (p16_and_64648_comb ^ p15_add_64534 & p15_add_64288 ^ p15_and_64529);
  assign p16_add_64629_comb = {p16_add_64607_comb[5:0] ^ p16_add_64607_comb[10:5] ^ p16_add_64607_comb[24:19], p16_add_64607_comb[31:27] ^ p16_add_64607_comb[4:0] ^ p16_add_64607_comb[18:14], p16_add_64607_comb[26:13] ^ p16_add_64607_comb[31:18] ^ p16_add_64607_comb[13:0], p16_add_64607_comb[12:6] ^ p16_add_64607_comb[17:11] ^ p16_add_64607_comb[31:25]} + (p16_add_64607_comb & p15_add_64487 ^ ~(p16_add_64607_comb | ~p15_add_64384));
  assign p16_add_64670_comb = p15_add_63831 + {p15_add_64552[16:7] ^ p15_add_64552[18:9], p15_add_64552[6:0] ^ p15_add_64552[8:2] ^ p15_add_64552[31:25], p15_add_64552[31:30] ^ p15_add_64552[1:0] ^ p15_add_64552[24:23], p15_add_64552[29:17] ^ p15_add_64552[31:19] ^ p15_add_64552[22:10]};
  assign p16_add_64653_comb = p15_add_64511 + p16_add_64652_comb;
  assign p16_add_64631_comb = p16_add_64629_comb + 32'h9bdc_06a7;
  assign p16_add_64671_comb = p15_add_63576 + p16_add_64670_comb;

  // Registers for pipe stage 16:
  reg [31:0] p16_add_64384;
  reg [31:0] p16_add_64487;
  reg [31:0] p16_add_64607;
  reg [31:0] p16_add_64512;
  reg [31:0] p16_add_64288;
  reg [31:0] p16_concat_63949;
  reg [31:0] p16_add_64430;
  reg [31:0] p16_add_64534;
  reg [31:0] p16_and_64648;
  reg [31:0] p16_add_64653;
  reg [1:0] p16_bit_slice_64535;
  reg [31:0] p16_add_64631;
  reg [31:0] p16_add_64325;
  reg [31:0] p16_add_64179;
  reg [31:0] p16_add_64162;
  reg [31:0] p16_add_64145;
  reg [31:0] p16_add_64128;
  reg [31:0] p16_add_64111;
  reg [31:0] p16_add_63848;
  reg [31:0] p16_add_64094;
  reg [31:0] p16_add_64671;
  reg [31:0] p16_add_64308;
  reg [31:0] p16_add_64552;
  reg [31:0] p16_add_64290;
  reg [31:0] p16_add_64289;
  reg [31:0] p16_add_64003;
  reg [31:0] p16_add_63985;
  reg [31:0] p16_add_63831;
  always_ff @ (posedge clk) begin
    p16_add_64384 <= p15_add_64384;
    p16_add_64487 <= p15_add_64487;
    p16_add_64607 <= p16_add_64607_comb;
    p16_add_64512 <= p15_add_64512;
    p16_add_64288 <= p15_add_64288;
    p16_concat_63949 <= p15_concat_63949;
    p16_add_64430 <= p15_add_64430;
    p16_add_64534 <= p15_add_64534;
    p16_and_64648 <= p16_and_64648_comb;
    p16_add_64653 <= p16_add_64653_comb;
    p16_bit_slice_64535 <= p15_bit_slice_64535;
    p16_add_64631 <= p16_add_64631_comb;
    p16_add_64325 <= p15_add_64325;
    p16_add_64179 <= p15_add_64179;
    p16_add_64162 <= p15_add_64162;
    p16_add_64145 <= p15_add_64145;
    p16_add_64128 <= p15_add_64128;
    p16_add_64111 <= p15_add_64111;
    p16_add_63848 <= p15_add_63848;
    p16_add_64094 <= p15_add_64094;
    p16_add_64671 <= p16_add_64671_comb;
    p16_add_64308 <= p15_add_64308;
    p16_add_64552 <= p15_add_64552;
    p16_add_64290 <= p15_add_64290;
    p16_add_64289 <= p15_add_64289;
    p16_add_64003 <= p15_add_64003;
    p16_add_63985 <= p15_add_63985;
    p16_add_63831 <= p15_add_63831;
  end

  // ===== Pipe stage 17:
  wire [31:0] p17_add_64728_comb;
  wire [31:0] p17_add_64729_comb;
  wire [31:0] p17_and_64770_comb;
  wire [31:0] p17_add_64774_comb;
  wire [31:0] p17_add_64792_comb;
  wire [31:0] p17_add_64753_comb;
  wire [31:0] p17_add_64775_comb;
  wire [31:0] p17_add_64810_comb;
  wire [31:0] p17_add_64793_comb;
  wire [31:0] p17_add_64751_comb;
  wire [31:0] p17_add_64752_comb;
  assign p17_add_64728_comb = p16_add_64631 + p16_add_64512;
  assign p17_add_64729_comb = p16_add_64288 + p17_add_64728_comb;
  assign p17_and_64770_comb = p16_add_64653 & p16_add_64534;
  assign p17_add_64774_comb = {p16_add_64653[1:0] ^ p16_add_64653[12:11] ^ p16_add_64653[21:20], p16_add_64653[31:21] ^ p16_add_64653[10:0] ^ p16_add_64653[19:9], p16_add_64653[20:12] ^ p16_add_64653[31:23] ^ p16_add_64653[8:0], p16_add_64653[11:2] ^ p16_add_64653[22:13] ^ p16_add_64653[31:22]} + (p17_and_64770_comb ^ p16_add_64653 & p16_add_64430 ^ p16_and_64648);
  assign p17_add_64792_comb = p16_add_64003 + {p16_add_64671[16:7] ^ p16_add_64671[18:9], p16_add_64671[6:0] ^ p16_add_64671[8:2] ^ p16_add_64671[31:25], p16_add_64671[31:30] ^ p16_add_64671[1:0] ^ p16_add_64671[24:23], p16_add_64671[29:17] ^ p16_add_64671[31:19] ^ p16_add_64671[22:10]};
  assign p17_add_64753_comb = p16_add_64487 + p16_add_63831;
  assign p17_add_64775_comb = p17_add_64728_comb + p17_add_64774_comb;
  assign p17_add_64810_comb = {p16_add_63985[6:4] ^ p16_add_63985[17:15], p16_add_63985[3:0] ^ p16_add_63985[14:11] ^ p16_add_63985[31:28], p16_add_63985[31:21] ^ p16_add_63985[10:0] ^ p16_add_63985[27:17], p16_add_63985[20:7] ^ p16_add_63985[31:18] ^ p16_add_63985[16:3]} + p16_add_63831;
  assign p17_add_64793_comb = p16_add_63848 + p17_add_64792_comb;
  assign p17_add_64751_comb = {p17_add_64729_comb[5:0] ^ p17_add_64729_comb[10:5] ^ p17_add_64729_comb[24:19], p17_add_64729_comb[31:27] ^ p17_add_64729_comb[4:0] ^ p17_add_64729_comb[18:14], p17_add_64729_comb[26:13] ^ p17_add_64729_comb[31:18] ^ p17_add_64729_comb[13:0], p17_add_64729_comb[12:6] ^ p17_add_64729_comb[17:11] ^ p17_add_64729_comb[31:25]} + p16_add_64384;
  assign p17_add_64752_comb = (p17_add_64729_comb & p16_add_64607 ^ ~(p17_add_64729_comb | ~p16_add_64487)) + p16_concat_63949;

  // Registers for pipe stage 17:
  reg [31:0] p17_add_64607;
  reg [31:0] p17_add_64729;
  reg [31:0] p17_add_64430;
  reg [31:0] p17_add_64753;
  reg [31:0] p17_add_64534;
  reg [31:0] p17_add_64653;
  reg [31:0] p17_and_64770;
  reg [31:0] p17_add_64775;
  reg [1:0] p17_bit_slice_64535;
  reg [31:0] p17_add_64810;
  reg [31:0] p17_add_64325;
  reg [31:0] p17_add_64179;
  reg [31:0] p17_add_64162;
  reg [31:0] p17_add_64145;
  reg [31:0] p17_add_64128;
  reg [31:0] p17_add_64111;
  reg [31:0] p17_add_64793;
  reg [31:0] p17_add_64094;
  reg [31:0] p17_add_64671;
  reg [31:0] p17_add_64308;
  reg [31:0] p17_add_64552;
  reg [31:0] p17_add_64290;
  reg [31:0] p17_add_64289;
  reg [31:0] p17_add_64003;
  reg [31:0] p17_add_63985;
  reg [31:0] p17_add_64751;
  reg [31:0] p17_add_64752;
  always_ff @ (posedge clk) begin
    p17_add_64607 <= p16_add_64607;
    p17_add_64729 <= p17_add_64729_comb;
    p17_add_64430 <= p16_add_64430;
    p17_add_64753 <= p17_add_64753_comb;
    p17_add_64534 <= p16_add_64534;
    p17_add_64653 <= p16_add_64653;
    p17_and_64770 <= p17_and_64770_comb;
    p17_add_64775 <= p17_add_64775_comb;
    p17_bit_slice_64535 <= p16_bit_slice_64535;
    p17_add_64810 <= p17_add_64810_comb;
    p17_add_64325 <= p16_add_64325;
    p17_add_64179 <= p16_add_64179;
    p17_add_64162 <= p16_add_64162;
    p17_add_64145 <= p16_add_64145;
    p17_add_64128 <= p16_add_64128;
    p17_add_64111 <= p16_add_64111;
    p17_add_64793 <= p17_add_64793_comb;
    p17_add_64094 <= p16_add_64094;
    p17_add_64671 <= p16_add_64671;
    p17_add_64308 <= p16_add_64308;
    p17_add_64552 <= p16_add_64552;
    p17_add_64290 <= p16_add_64290;
    p17_add_64289 <= p16_add_64289;
    p17_add_64003 <= p16_add_64003;
    p17_add_63985 <= p16_add_63985;
    p17_add_64751 <= p17_add_64751_comb;
    p17_add_64752 <= p17_add_64752_comb;
  end

  // ===== Pipe stage 18:
  wire [31:0] p18_add_64865_comb;
  wire [31:0] p18_add_64866_comb;
  wire [31:0] p18_and_64905_comb;
  wire [31:0] p18_add_64909_comb;
  wire [31:0] p18_add_64927_comb;
  wire [31:0] p18_add_64888_comb;
  wire [31:0] p18_add_64910_comb;
  wire [31:0] p18_add_64928_comb;
  assign p18_add_64865_comb = p17_add_64751 + p17_add_64752;
  assign p18_add_64866_comb = p17_add_64430 + p18_add_64865_comb;
  assign p18_and_64905_comb = p17_add_64775 & p17_add_64653;
  assign p18_add_64909_comb = {p17_add_64775[1:0] ^ p17_add_64775[12:11] ^ p17_add_64775[21:20], p17_add_64775[31:21] ^ p17_add_64775[10:0] ^ p17_add_64775[19:9], p17_add_64775[20:12] ^ p17_add_64775[31:23] ^ p17_add_64775[8:0], p17_add_64775[11:2] ^ p17_add_64775[22:13] ^ p17_add_64775[31:22]} + (p18_and_64905_comb ^ p17_add_64775 & p17_add_64534 ^ p17_and_64770);
  assign p18_add_64927_comb = p17_add_64290 + {p17_add_64793[16:7] ^ p17_add_64793[18:9], p17_add_64793[6:0] ^ p17_add_64793[8:2] ^ p17_add_64793[31:25], p17_add_64793[31:30] ^ p17_add_64793[1:0] ^ p17_add_64793[24:23], p17_add_64793[29:17] ^ p17_add_64793[31:19] ^ p17_add_64793[22:10]};
  assign p18_add_64888_comb = {p18_add_64866_comb[5:0] ^ p18_add_64866_comb[10:5] ^ p18_add_64866_comb[24:19], p18_add_64866_comb[31:27] ^ p18_add_64866_comb[4:0] ^ p18_add_64866_comb[18:14], p18_add_64866_comb[26:13] ^ p18_add_64866_comb[31:18] ^ p18_add_64866_comb[13:0], p18_add_64866_comb[12:6] ^ p18_add_64866_comb[17:11] ^ p18_add_64866_comb[31:25]} + (p18_add_64866_comb & p17_add_64729 ^ ~(p18_add_64866_comb | ~p17_add_64607));
  assign p18_add_64910_comb = p18_add_64865_comb + p18_add_64909_comb;
  assign p18_add_64928_comb = p17_add_64128 + p18_add_64927_comb;

  // Registers for pipe stage 18:
  reg [31:0] p18_add_64607;
  reg [31:0] p18_add_64729;
  reg [31:0] p18_add_64866;
  reg [31:0] p18_add_64888;
  reg [31:0] p18_add_64753;
  reg [31:0] p18_add_64534;
  reg [31:0] p18_add_64653;
  reg [31:0] p18_add_64775;
  reg [1:0] p18_bit_slice_64535;
  reg [31:0] p18_and_64905;
  reg [31:0] p18_add_64910;
  reg [31:0] p18_add_64810;
  reg [31:0] p18_add_64325;
  reg [31:0] p18_add_64179;
  reg [31:0] p18_add_64162;
  reg [31:0] p18_add_64145;
  reg [31:0] p18_add_64928;
  reg [31:0] p18_add_64111;
  reg [31:0] p18_add_64793;
  reg [31:0] p18_add_64094;
  reg [31:0] p18_add_64671;
  reg [31:0] p18_add_64308;
  reg [31:0] p18_add_64552;
  reg [31:0] p18_add_64290;
  reg [31:0] p18_add_64289;
  reg [31:0] p18_add_64003;
  reg [31:0] p18_add_63985;
  always_ff @ (posedge clk) begin
    p18_add_64607 <= p17_add_64607;
    p18_add_64729 <= p17_add_64729;
    p18_add_64866 <= p18_add_64866_comb;
    p18_add_64888 <= p18_add_64888_comb;
    p18_add_64753 <= p17_add_64753;
    p18_add_64534 <= p17_add_64534;
    p18_add_64653 <= p17_add_64653;
    p18_add_64775 <= p17_add_64775;
    p18_bit_slice_64535 <= p17_bit_slice_64535;
    p18_and_64905 <= p18_and_64905_comb;
    p18_add_64910 <= p18_add_64910_comb;
    p18_add_64810 <= p17_add_64810;
    p18_add_64325 <= p17_add_64325;
    p18_add_64179 <= p17_add_64179;
    p18_add_64162 <= p17_add_64162;
    p18_add_64145 <= p17_add_64145;
    p18_add_64928 <= p18_add_64928_comb;
    p18_add_64111 <= p17_add_64111;
    p18_add_64793 <= p17_add_64793;
    p18_add_64094 <= p17_add_64094;
    p18_add_64671 <= p17_add_64671;
    p18_add_64308 <= p17_add_64308;
    p18_add_64552 <= p17_add_64552;
    p18_add_64290 <= p17_add_64290;
    p18_add_64289 <= p17_add_64289;
    p18_add_64003 <= p17_add_64003;
    p18_add_63985 <= p17_add_63985;
  end

  // ===== Pipe stage 19:
  wire [31:0] p19_and_65006_comb;
  wire [31:0] p19_add_64984_comb;
  wire [31:0] p19_add_64985_comb;
  wire [31:0] p19_add_65010_comb;
  wire [31:0] p19_add_65028_comb;
  wire [31:0] p19_add_64986_comb;
  wire [30:0] p19_add_64989_comb;
  wire [31:0] p19_add_65011_comb;
  wire [31:0] p19_add_65029_comb;
  assign p19_and_65006_comb = p18_add_64910 & p18_add_64775;
  assign p19_add_64984_comb = p18_add_64888 + 32'he49b_69c1;
  assign p19_add_64985_comb = p19_add_64984_comb + p18_add_64753;
  assign p19_add_65010_comb = {p18_add_64910[1:0] ^ p18_add_64910[12:11] ^ p18_add_64910[21:20], p18_add_64910[31:21] ^ p18_add_64910[10:0] ^ p18_add_64910[19:9], p18_add_64910[20:12] ^ p18_add_64910[31:23] ^ p18_add_64910[8:0], p18_add_64910[11:2] ^ p18_add_64910[22:13] ^ p18_add_64910[31:22]} + (p19_and_65006_comb ^ p18_add_64910 & p18_add_64653 ^ p18_and_64905);
  assign p19_add_65028_comb = p18_add_64308 + {p18_add_64928[16:7] ^ p18_add_64928[18:9], p18_add_64928[6:0] ^ p18_add_64928[8:2] ^ p18_add_64928[31:25], p18_add_64928[31:30] ^ p18_add_64928[1:0] ^ p18_add_64928[24:23], p18_add_64928[29:17] ^ p18_add_64928[31:19] ^ p18_add_64928[22:10]};
  assign p19_add_64986_comb = p18_add_64534 + p19_add_64985_comb;
  assign p19_add_64989_comb = p18_add_63985[31:1] + 31'h77df_23c3;
  assign p19_add_65011_comb = p19_add_64985_comb + p19_add_65010_comb;
  assign p19_add_65029_comb = p18_add_64162 + p19_add_65028_comb;

  // Registers for pipe stage 19:
  reg [31:0] p19_add_64607;
  reg [31:0] p19_add_64729;
  reg [31:0] p19_add_64866;
  reg [31:0] p19_add_64986;
  reg [30:0] p19_add_64989;
  reg [31:0] p19_add_64653;
  reg [31:0] p19_add_64775;
  reg [1:0] p19_bit_slice_64535;
  reg [31:0] p19_add_64910;
  reg [31:0] p19_and_65006;
  reg [31:0] p19_add_65011;
  reg [31:0] p19_add_64810;
  reg [31:0] p19_add_64325;
  reg [31:0] p19_add_64179;
  reg [31:0] p19_add_65029;
  reg [31:0] p19_add_64145;
  reg [31:0] p19_add_64928;
  reg [31:0] p19_add_64111;
  reg [31:0] p19_add_64793;
  reg [31:0] p19_add_64094;
  reg [31:0] p19_add_64671;
  reg [31:0] p19_add_64308;
  reg [31:0] p19_add_64552;
  reg [31:0] p19_add_64290;
  reg [31:0] p19_add_64289;
  reg [31:0] p19_add_64003;
  reg [31:0] p19_add_63985;
  always_ff @ (posedge clk) begin
    p19_add_64607 <= p18_add_64607;
    p19_add_64729 <= p18_add_64729;
    p19_add_64866 <= p18_add_64866;
    p19_add_64986 <= p19_add_64986_comb;
    p19_add_64989 <= p19_add_64989_comb;
    p19_add_64653 <= p18_add_64653;
    p19_add_64775 <= p18_add_64775;
    p19_bit_slice_64535 <= p18_bit_slice_64535;
    p19_add_64910 <= p18_add_64910;
    p19_and_65006 <= p19_and_65006_comb;
    p19_add_65011 <= p19_add_65011_comb;
    p19_add_64810 <= p18_add_64810;
    p19_add_64325 <= p18_add_64325;
    p19_add_64179 <= p18_add_64179;
    p19_add_65029 <= p19_add_65029_comb;
    p19_add_64145 <= p18_add_64145;
    p19_add_64928 <= p18_add_64928;
    p19_add_64111 <= p18_add_64111;
    p19_add_64793 <= p18_add_64793;
    p19_add_64094 <= p18_add_64094;
    p19_add_64671 <= p18_add_64671;
    p19_add_64308 <= p18_add_64308;
    p19_add_64552 <= p18_add_64552;
    p19_add_64290 <= p18_add_64290;
    p19_add_64289 <= p18_add_64289;
    p19_add_64003 <= p18_add_64003;
    p19_add_63985 <= p18_add_63985;
  end

  // ===== Pipe stage 20:
  wire [31:0] p20_and_65130_comb;
  wire [31:0] p20_add_65107_comb;
  wire [31:0] p20_add_65108_comb;
  wire [31:0] p20_add_65109_comb;
  wire [31:0] p20_add_65134_comb;
  wire [31:0] p20_add_65110_comb;
  wire [30:0] p20_add_65113_comb;
  wire [31:0] p20_add_65135_comb;
  assign p20_and_65130_comb = p19_add_65011 & p19_add_64910;
  assign p20_add_65107_comb = {p19_add_64986[5:0] ^ p19_add_64986[10:5] ^ p19_add_64986[24:19], p19_add_64986[31:27] ^ p19_add_64986[4:0] ^ p19_add_64986[18:14], p19_add_64986[26:13] ^ p19_add_64986[31:18] ^ p19_add_64986[13:0], p19_add_64986[12:6] ^ p19_add_64986[17:11] ^ p19_add_64986[31:25]} + p19_add_64607;
  assign p20_add_65108_comb = (p19_add_64986 & p19_add_64866 ^ ~(p19_add_64986 | ~p19_add_64729)) + {p19_add_64989, p19_add_63985[0]};
  assign p20_add_65109_comb = p20_add_65107_comb + p20_add_65108_comb;
  assign p20_add_65134_comb = {p19_add_65011[1:0] ^ p19_add_65011[12:11] ^ p19_add_65011[21:20], p19_add_65011[31:21] ^ p19_add_65011[10:0] ^ p19_add_65011[19:9], p19_add_65011[20:12] ^ p19_add_65011[31:23] ^ p19_add_65011[8:0], p19_add_65011[11:2] ^ p19_add_65011[22:13] ^ p19_add_65011[31:22]} + (p20_and_65130_comb ^ p19_add_65011 & p19_add_64775 ^ p19_and_65006);
  assign p20_add_65110_comb = p19_add_64653 + p20_add_65109_comb;
  assign p20_add_65113_comb = p19_add_64003[31:1] + 31'h07e0_cee3;
  assign p20_add_65135_comb = p20_add_65109_comb + p20_add_65134_comb;

  // Registers for pipe stage 20:
  reg [31:0] p20_add_64729;
  reg [31:0] p20_add_64866;
  reg [31:0] p20_add_64986;
  reg [31:0] p20_add_65110;
  reg [30:0] p20_add_65113;
  reg [31:0] p20_add_64775;
  reg [1:0] p20_bit_slice_64535;
  reg [31:0] p20_add_64910;
  reg [31:0] p20_add_65011;
  reg [31:0] p20_and_65130;
  reg [31:0] p20_add_65135;
  reg [31:0] p20_add_64810;
  reg [31:0] p20_add_64325;
  reg [31:0] p20_add_64179;
  reg [31:0] p20_add_65029;
  reg [31:0] p20_add_64145;
  reg [31:0] p20_add_64928;
  reg [31:0] p20_add_64111;
  reg [31:0] p20_add_64793;
  reg [31:0] p20_add_64094;
  reg [31:0] p20_add_64671;
  reg [31:0] p20_add_64308;
  reg [31:0] p20_add_64552;
  reg [31:0] p20_add_64290;
  reg [31:0] p20_add_64289;
  reg [31:0] p20_add_64003;
  reg [31:0] p20_add_63985;
  always_ff @ (posedge clk) begin
    p20_add_64729 <= p19_add_64729;
    p20_add_64866 <= p19_add_64866;
    p20_add_64986 <= p19_add_64986;
    p20_add_65110 <= p20_add_65110_comb;
    p20_add_65113 <= p20_add_65113_comb;
    p20_add_64775 <= p19_add_64775;
    p20_bit_slice_64535 <= p19_bit_slice_64535;
    p20_add_64910 <= p19_add_64910;
    p20_add_65011 <= p19_add_65011;
    p20_and_65130 <= p20_and_65130_comb;
    p20_add_65135 <= p20_add_65135_comb;
    p20_add_64810 <= p19_add_64810;
    p20_add_64325 <= p19_add_64325;
    p20_add_64179 <= p19_add_64179;
    p20_add_65029 <= p19_add_65029;
    p20_add_64145 <= p19_add_64145;
    p20_add_64928 <= p19_add_64928;
    p20_add_64111 <= p19_add_64111;
    p20_add_64793 <= p19_add_64793;
    p20_add_64094 <= p19_add_64094;
    p20_add_64671 <= p19_add_64671;
    p20_add_64308 <= p19_add_64308;
    p20_add_64552 <= p19_add_64552;
    p20_add_64290 <= p19_add_64290;
    p20_add_64289 <= p19_add_64289;
    p20_add_64003 <= p19_add_64003;
    p20_add_63985 <= p19_add_63985;
  end

  // ===== Pipe stage 21:
  wire [31:0] p21_and_65237_comb;
  wire [31:0] p21_add_65213_comb;
  wire [31:0] p21_add_65214_comb;
  wire [31:0] p21_add_65215_comb;
  wire [29:0] p21_add_65219_comb;
  wire [31:0] p21_add_65241_comb;
  wire [31:0] p21_add_65216_comb;
  wire [31:0] p21_concat_65220_comb;
  wire [31:0] p21_add_65242_comb;
  assign p21_and_65237_comb = p20_add_65135 & p20_add_65011;
  assign p21_add_65213_comb = {p20_add_65110[5:0] ^ p20_add_65110[10:5] ^ p20_add_65110[24:19], p20_add_65110[31:27] ^ p20_add_65110[4:0] ^ p20_add_65110[18:14], p20_add_65110[26:13] ^ p20_add_65110[31:18] ^ p20_add_65110[13:0], p20_add_65110[12:6] ^ p20_add_65110[17:11] ^ p20_add_65110[31:25]} + p20_add_64729;
  assign p21_add_65214_comb = (p20_add_65110 & p20_add_64986 ^ ~(p20_add_65110 | ~p20_add_64866)) + {p20_add_65113, p20_add_64003[0]};
  assign p21_add_65215_comb = p21_add_65213_comb + p21_add_65214_comb;
  assign p21_add_65219_comb = p20_add_64289[31:2] + 30'h0903_2873;
  assign p21_add_65241_comb = {p20_add_65135[1:0] ^ p20_add_65135[12:11] ^ p20_add_65135[21:20], p20_add_65135[31:21] ^ p20_add_65135[10:0] ^ p20_add_65135[19:9], p20_add_65135[20:12] ^ p20_add_65135[31:23] ^ p20_add_65135[8:0], p20_add_65135[11:2] ^ p20_add_65135[22:13] ^ p20_add_65135[31:22]} + (p21_and_65237_comb ^ p20_add_65135 & p20_add_64910 ^ p20_and_65130);
  assign p21_add_65216_comb = p20_add_64775 + p21_add_65215_comb;
  assign p21_concat_65220_comb = {p21_add_65219_comb, p20_bit_slice_64535};
  assign p21_add_65242_comb = p21_add_65215_comb + p21_add_65241_comb;

  // Registers for pipe stage 21:
  reg [31:0] p21_add_64866;
  reg [31:0] p21_add_64986;
  reg [31:0] p21_add_65110;
  reg [31:0] p21_add_65216;
  reg [31:0] p21_concat_65220;
  reg [31:0] p21_add_64910;
  reg [31:0] p21_add_65011;
  reg [31:0] p21_add_65135;
  reg [31:0] p21_and_65237;
  reg [31:0] p21_add_65242;
  reg [31:0] p21_add_64810;
  reg [31:0] p21_add_64325;
  reg [31:0] p21_add_64179;
  reg [31:0] p21_add_65029;
  reg [31:0] p21_add_64145;
  reg [31:0] p21_add_64928;
  reg [31:0] p21_add_64111;
  reg [31:0] p21_add_64793;
  reg [31:0] p21_add_64094;
  reg [31:0] p21_add_64671;
  reg [31:0] p21_add_64308;
  reg [31:0] p21_add_64552;
  reg [31:0] p21_add_64290;
  reg [31:0] p21_add_64289;
  reg [31:0] p21_add_64003;
  reg [31:0] p21_add_63985;
  always_ff @ (posedge clk) begin
    p21_add_64866 <= p20_add_64866;
    p21_add_64986 <= p20_add_64986;
    p21_add_65110 <= p20_add_65110;
    p21_add_65216 <= p21_add_65216_comb;
    p21_concat_65220 <= p21_concat_65220_comb;
    p21_add_64910 <= p20_add_64910;
    p21_add_65011 <= p20_add_65011;
    p21_add_65135 <= p20_add_65135;
    p21_and_65237 <= p21_and_65237_comb;
    p21_add_65242 <= p21_add_65242_comb;
    p21_add_64810 <= p20_add_64810;
    p21_add_64325 <= p20_add_64325;
    p21_add_64179 <= p20_add_64179;
    p21_add_65029 <= p20_add_65029;
    p21_add_64145 <= p20_add_64145;
    p21_add_64928 <= p20_add_64928;
    p21_add_64111 <= p20_add_64111;
    p21_add_64793 <= p20_add_64793;
    p21_add_64094 <= p20_add_64094;
    p21_add_64671 <= p20_add_64671;
    p21_add_64308 <= p20_add_64308;
    p21_add_64552 <= p20_add_64552;
    p21_add_64290 <= p20_add_64290;
    p21_add_64289 <= p20_add_64289;
    p21_add_64003 <= p20_add_64003;
    p21_add_63985 <= p20_add_63985;
  end

  // ===== Pipe stage 22:
  wire [31:0] p22_and_65337_comb;
  wire [31:0] p22_add_65316_comb;
  wire [31:0] p22_add_65317_comb;
  wire [31:0] p22_add_65318_comb;
  wire [31:0] p22_add_65341_comb;
  wire [31:0] p22_add_65319_comb;
  wire [31:0] p22_add_65320_comb;
  wire [31:0] p22_add_65342_comb;
  assign p22_and_65337_comb = p21_add_65242 & p21_add_65135;
  assign p22_add_65316_comb = {p21_add_65216[5:0] ^ p21_add_65216[10:5] ^ p21_add_65216[24:19], p21_add_65216[31:27] ^ p21_add_65216[4:0] ^ p21_add_65216[18:14], p21_add_65216[26:13] ^ p21_add_65216[31:18] ^ p21_add_65216[13:0], p21_add_65216[12:6] ^ p21_add_65216[17:11] ^ p21_add_65216[31:25]} + p21_add_64866;
  assign p22_add_65317_comb = (p21_add_65216 & p21_add_65110 ^ ~(p21_add_65216 | ~p21_add_64986)) + p21_concat_65220;
  assign p22_add_65318_comb = p22_add_65316_comb + p22_add_65317_comb;
  assign p22_add_65341_comb = {p21_add_65242[1:0] ^ p21_add_65242[12:11] ^ p21_add_65242[21:20], p21_add_65242[31:21] ^ p21_add_65242[10:0] ^ p21_add_65242[19:9], p21_add_65242[20:12] ^ p21_add_65242[31:23] ^ p21_add_65242[8:0], p21_add_65242[11:2] ^ p21_add_65242[22:13] ^ p21_add_65242[31:22]} + (p22_and_65337_comb ^ p21_add_65242 & p21_add_65011 ^ p21_and_65237);
  assign p22_add_65319_comb = p21_add_64910 + p22_add_65318_comb;
  assign p22_add_65320_comb = p21_add_64986 + p21_add_64290;
  assign p22_add_65342_comb = p22_add_65318_comb + p22_add_65341_comb;

  // Registers for pipe stage 22:
  reg [31:0] p22_add_65110;
  reg [31:0] p22_add_65216;
  reg [31:0] p22_add_65319;
  reg [31:0] p22_add_65320;
  reg [31:0] p22_add_65011;
  reg [31:0] p22_add_65135;
  reg [31:0] p22_add_65242;
  reg [31:0] p22_and_65337;
  reg [31:0] p22_add_65342;
  reg [31:0] p22_add_64810;
  reg [31:0] p22_add_64325;
  reg [31:0] p22_add_64179;
  reg [31:0] p22_add_65029;
  reg [31:0] p22_add_64145;
  reg [31:0] p22_add_64928;
  reg [31:0] p22_add_64111;
  reg [31:0] p22_add_64793;
  reg [31:0] p22_add_64094;
  reg [31:0] p22_add_64671;
  reg [31:0] p22_add_64308;
  reg [31:0] p22_add_64552;
  reg [31:0] p22_add_64290;
  reg [31:0] p22_add_64289;
  reg [31:0] p22_add_64003;
  reg [31:0] p22_add_63985;
  always_ff @ (posedge clk) begin
    p22_add_65110 <= p21_add_65110;
    p22_add_65216 <= p21_add_65216;
    p22_add_65319 <= p22_add_65319_comb;
    p22_add_65320 <= p22_add_65320_comb;
    p22_add_65011 <= p21_add_65011;
    p22_add_65135 <= p21_add_65135;
    p22_add_65242 <= p21_add_65242;
    p22_and_65337 <= p22_and_65337_comb;
    p22_add_65342 <= p22_add_65342_comb;
    p22_add_64810 <= p21_add_64810;
    p22_add_64325 <= p21_add_64325;
    p22_add_64179 <= p21_add_64179;
    p22_add_65029 <= p21_add_65029;
    p22_add_64145 <= p21_add_64145;
    p22_add_64928 <= p21_add_64928;
    p22_add_64111 <= p21_add_64111;
    p22_add_64793 <= p21_add_64793;
    p22_add_64094 <= p21_add_64094;
    p22_add_64671 <= p21_add_64671;
    p22_add_64308 <= p21_add_64308;
    p22_add_64552 <= p21_add_64552;
    p22_add_64290 <= p21_add_64290;
    p22_add_64289 <= p21_add_64289;
    p22_add_64003 <= p21_add_64003;
    p22_add_63985 <= p21_add_63985;
  end

  // ===== Pipe stage 23:
  wire [31:0] p23_add_65414_comb;
  wire [31:0] p23_add_65416_comb;
  wire [31:0] p23_add_65417_comb;
  assign p23_add_65414_comb = {p22_add_65319[5:0] ^ p22_add_65319[10:5] ^ p22_add_65319[24:19], p22_add_65319[31:27] ^ p22_add_65319[4:0] ^ p22_add_65319[18:14], p22_add_65319[26:13] ^ p22_add_65319[31:18] ^ p22_add_65319[13:0], p22_add_65319[12:6] ^ p22_add_65319[17:11] ^ p22_add_65319[31:25]} + (p22_add_65319 & p22_add_65216 ^ ~(p22_add_65319 | ~p22_add_65110));
  assign p23_add_65416_comb = p23_add_65414_comb + 32'h2de9_2c6f;
  assign p23_add_65417_comb = p23_add_65416_comb + p22_add_65320;

  // Registers for pipe stage 23:
  reg [31:0] p23_add_65110;
  reg [31:0] p23_add_65216;
  reg [31:0] p23_add_65319;
  reg [31:0] p23_add_65011;
  reg [31:0] p23_add_65417;
  reg [31:0] p23_add_65135;
  reg [31:0] p23_add_65242;
  reg [31:0] p23_and_65337;
  reg [31:0] p23_add_65342;
  reg [31:0] p23_add_64810;
  reg [31:0] p23_add_64325;
  reg [31:0] p23_add_64179;
  reg [31:0] p23_add_65029;
  reg [31:0] p23_add_64145;
  reg [31:0] p23_add_64928;
  reg [31:0] p23_add_64111;
  reg [31:0] p23_add_64793;
  reg [31:0] p23_add_64094;
  reg [31:0] p23_add_64671;
  reg [31:0] p23_add_64308;
  reg [31:0] p23_add_64552;
  reg [31:0] p23_add_64290;
  reg [31:0] p23_add_64289;
  reg [31:0] p23_add_64003;
  reg [31:0] p23_add_63985;
  always_ff @ (posedge clk) begin
    p23_add_65110 <= p22_add_65110;
    p23_add_65216 <= p22_add_65216;
    p23_add_65319 <= p22_add_65319;
    p23_add_65011 <= p22_add_65011;
    p23_add_65417 <= p23_add_65417_comb;
    p23_add_65135 <= p22_add_65135;
    p23_add_65242 <= p22_add_65242;
    p23_and_65337 <= p22_and_65337;
    p23_add_65342 <= p22_add_65342;
    p23_add_64810 <= p22_add_64810;
    p23_add_64325 <= p22_add_64325;
    p23_add_64179 <= p22_add_64179;
    p23_add_65029 <= p22_add_65029;
    p23_add_64145 <= p22_add_64145;
    p23_add_64928 <= p22_add_64928;
    p23_add_64111 <= p22_add_64111;
    p23_add_64793 <= p22_add_64793;
    p23_add_64094 <= p22_add_64094;
    p23_add_64671 <= p22_add_64671;
    p23_add_64308 <= p22_add_64308;
    p23_add_64552 <= p22_add_64552;
    p23_add_64290 <= p22_add_64290;
    p23_add_64289 <= p22_add_64289;
    p23_add_64003 <= p22_add_64003;
    p23_add_63985 <= p22_add_63985;
  end

  // ===== Pipe stage 24:
  wire [31:0] p24_add_65468_comb;
  wire [31:0] p24_and_65514_comb;
  wire [30:0] p24_add_65490_comb;
  wire [31:0] p24_add_65518_comb;
  wire [31:0] p24_add_65495_comb;
  wire [31:0] p24_add_65496_comb;
  wire [31:0] p24_add_65519_comb;
  wire [31:0] p24_add_65497_comb;
  assign p24_add_65468_comb = p23_add_65011 + p23_add_65417;
  assign p24_and_65514_comb = p23_add_65342 & p23_add_65242;
  assign p24_add_65490_comb = p23_add_64552[31:1] + 31'h253a_4255;
  assign p24_add_65518_comb = {p23_add_65342[1:0] ^ p23_add_65342[12:11] ^ p23_add_65342[21:20], p23_add_65342[31:21] ^ p23_add_65342[10:0] ^ p23_add_65342[19:9], p23_add_65342[20:12] ^ p23_add_65342[31:23] ^ p23_add_65342[8:0], p23_add_65342[11:2] ^ p23_add_65342[22:13] ^ p23_add_65342[31:22]} + (p24_and_65514_comb ^ p23_add_65342 & p23_add_65135 ^ p23_and_65337);
  assign p24_add_65495_comb = {p24_add_65468_comb[5:0] ^ p24_add_65468_comb[10:5] ^ p24_add_65468_comb[24:19], p24_add_65468_comb[31:27] ^ p24_add_65468_comb[4:0] ^ p24_add_65468_comb[18:14], p24_add_65468_comb[26:13] ^ p24_add_65468_comb[31:18] ^ p24_add_65468_comb[13:0], p24_add_65468_comb[12:6] ^ p24_add_65468_comb[17:11] ^ p24_add_65468_comb[31:25]} + p23_add_65110;
  assign p24_add_65496_comb = (p24_add_65468_comb & p23_add_65319 ^ ~(p24_add_65468_comb | ~p23_add_65216)) + {p24_add_65490_comb, p23_add_64552[0]};
  assign p24_add_65519_comb = p23_add_65417 + p24_add_65518_comb;
  assign p24_add_65497_comb = p24_add_65495_comb + p24_add_65496_comb;

  // Registers for pipe stage 24:
  reg [31:0] p24_add_65216;
  reg [31:0] p24_add_65319;
  reg [31:0] p24_add_65468;
  reg [31:0] p24_add_65135;
  reg [31:0] p24_add_65242;
  reg [31:0] p24_add_65342;
  reg [31:0] p24_and_65514;
  reg [31:0] p24_add_65519;
  reg [31:0] p24_add_64810;
  reg [31:0] p24_add_64325;
  reg [31:0] p24_add_64179;
  reg [31:0] p24_add_65029;
  reg [31:0] p24_add_64145;
  reg [31:0] p24_add_64928;
  reg [31:0] p24_add_64111;
  reg [31:0] p24_add_64793;
  reg [31:0] p24_add_64094;
  reg [31:0] p24_add_64671;
  reg [31:0] p24_add_64308;
  reg [31:0] p24_add_65497;
  reg [31:0] p24_add_64552;
  reg [31:0] p24_add_64290;
  reg [31:0] p24_add_64289;
  reg [31:0] p24_add_64003;
  reg [31:0] p24_add_63985;
  always_ff @ (posedge clk) begin
    p24_add_65216 <= p23_add_65216;
    p24_add_65319 <= p23_add_65319;
    p24_add_65468 <= p24_add_65468_comb;
    p24_add_65135 <= p23_add_65135;
    p24_add_65242 <= p23_add_65242;
    p24_add_65342 <= p23_add_65342;
    p24_and_65514 <= p24_and_65514_comb;
    p24_add_65519 <= p24_add_65519_comb;
    p24_add_64810 <= p23_add_64810;
    p24_add_64325 <= p23_add_64325;
    p24_add_64179 <= p23_add_64179;
    p24_add_65029 <= p23_add_65029;
    p24_add_64145 <= p23_add_64145;
    p24_add_64928 <= p23_add_64928;
    p24_add_64111 <= p23_add_64111;
    p24_add_64793 <= p23_add_64793;
    p24_add_64094 <= p23_add_64094;
    p24_add_64671 <= p23_add_64671;
    p24_add_64308 <= p23_add_64308;
    p24_add_65497 <= p24_add_65497_comb;
    p24_add_64552 <= p23_add_64552;
    p24_add_64290 <= p23_add_64290;
    p24_add_64289 <= p23_add_64289;
    p24_add_64003 <= p23_add_64003;
    p24_add_63985 <= p23_add_63985;
  end

  // ===== Pipe stage 25:
  wire [31:0] p25_add_65570_comb;
  wire [31:0] p25_and_65633_comb;
  wire [29:0] p25_add_65592_comb;
  wire [31:0] p25_add_65637_comb;
  wire [31:0] p25_add_65615_comb;
  wire [31:0] p25_add_65597_comb;
  wire [31:0] p25_add_65598_comb;
  wire [31:0] p25_add_65638_comb;
  wire [31:0] p25_add_65672_comb;
  wire [31:0] p25_add_65655_comb;
  wire [31:0] p25_add_65616_comb;
  wire [31:0] p25_add_65599_comb;
  assign p25_add_65570_comb = p24_add_65135 + p24_add_65497;
  assign p25_and_65633_comb = p24_add_65519 & p24_add_65342;
  assign p25_add_65592_comb = p24_add_64308[31:2] + 30'h172c_2a77;
  assign p25_add_65637_comb = {p24_add_65519[1:0] ^ p24_add_65519[12:11] ^ p24_add_65519[21:20], p24_add_65519[31:21] ^ p24_add_65519[10:0] ^ p24_add_65519[19:9], p24_add_65519[20:12] ^ p24_add_65519[31:23] ^ p24_add_65519[8:0], p24_add_65519[11:2] ^ p24_add_65519[22:13] ^ p24_add_65519[31:22]} + (p25_and_65633_comb ^ p24_add_65519 & p24_add_65242 ^ p24_and_65514);
  assign p25_add_65615_comb = p24_add_63985 + {p24_add_64308[16:7] ^ p24_add_64308[18:9], p24_add_64308[6:0] ^ p24_add_64308[8:2] ^ p24_add_64308[31:25], p24_add_64308[31:30] ^ p24_add_64308[1:0] ^ p24_add_64308[24:23], p24_add_64308[29:17] ^ p24_add_64308[31:19] ^ p24_add_64308[22:10]};
  assign p25_add_65597_comb = {p25_add_65570_comb[5:0] ^ p25_add_65570_comb[10:5] ^ p25_add_65570_comb[24:19], p25_add_65570_comb[31:27] ^ p25_add_65570_comb[4:0] ^ p25_add_65570_comb[18:14], p25_add_65570_comb[26:13] ^ p25_add_65570_comb[31:18] ^ p25_add_65570_comb[13:0], p25_add_65570_comb[12:6] ^ p25_add_65570_comb[17:11] ^ p25_add_65570_comb[31:25]} + p24_add_65216;
  assign p25_add_65598_comb = (p25_add_65570_comb & p24_add_65468 ^ ~(p25_add_65570_comb | ~p24_add_65319)) + {p25_add_65592_comb, p24_add_64308[1:0]};
  assign p25_add_65638_comb = p24_add_65497 + p25_add_65637_comb;
  assign p25_add_65672_comb = {p24_add_64289[6:4] ^ p24_add_64289[17:15], p24_add_64289[3:0] ^ p24_add_64289[14:11] ^ p24_add_64289[31:28], p24_add_64289[31:21] ^ p24_add_64289[10:0] ^ p24_add_64289[27:17], p24_add_64289[20:7] ^ p24_add_64289[31:18] ^ p24_add_64289[16:3]} + p24_add_64003;
  assign p25_add_65655_comb = {p24_add_64003[6:4] ^ p24_add_64003[17:15], p24_add_64003[3:0] ^ p24_add_64003[14:11] ^ p24_add_64003[31:28], p24_add_64003[31:21] ^ p24_add_64003[10:0] ^ p24_add_64003[27:17], p24_add_64003[20:7] ^ p24_add_64003[31:18] ^ p24_add_64003[16:3]} + p24_add_63985;
  assign p25_add_65616_comb = p24_add_64094 + p25_add_65615_comb;
  assign p25_add_65599_comb = p25_add_65597_comb + p25_add_65598_comb;

  // Registers for pipe stage 25:
  reg [31:0] p25_add_65319;
  reg [31:0] p25_add_65468;
  reg [31:0] p25_add_65570;
  reg [31:0] p25_add_65242;
  reg [31:0] p25_add_65342;
  reg [31:0] p25_add_65519;
  reg [31:0] p25_and_65633;
  reg [31:0] p25_add_65638;
  reg [31:0] p25_add_65672;
  reg [31:0] p25_add_65655;
  reg [31:0] p25_add_64810;
  reg [31:0] p25_add_64325;
  reg [31:0] p25_add_64179;
  reg [31:0] p25_add_65029;
  reg [31:0] p25_add_64145;
  reg [31:0] p25_add_64928;
  reg [31:0] p25_add_64111;
  reg [31:0] p25_add_64793;
  reg [31:0] p25_add_65616;
  reg [31:0] p25_add_64671;
  reg [31:0] p25_add_65599;
  reg [31:0] p25_add_64308;
  reg [31:0] p25_add_64552;
  reg [31:0] p25_add_64290;
  reg [31:0] p25_add_64289;
  always_ff @ (posedge clk) begin
    p25_add_65319 <= p24_add_65319;
    p25_add_65468 <= p24_add_65468;
    p25_add_65570 <= p25_add_65570_comb;
    p25_add_65242 <= p24_add_65242;
    p25_add_65342 <= p24_add_65342;
    p25_add_65519 <= p24_add_65519;
    p25_and_65633 <= p25_and_65633_comb;
    p25_add_65638 <= p25_add_65638_comb;
    p25_add_65672 <= p25_add_65672_comb;
    p25_add_65655 <= p25_add_65655_comb;
    p25_add_64810 <= p24_add_64810;
    p25_add_64325 <= p24_add_64325;
    p25_add_64179 <= p24_add_64179;
    p25_add_65029 <= p24_add_65029;
    p25_add_64145 <= p24_add_64145;
    p25_add_64928 <= p24_add_64928;
    p25_add_64111 <= p24_add_64111;
    p25_add_64793 <= p24_add_64793;
    p25_add_65616 <= p25_add_65616_comb;
    p25_add_64671 <= p24_add_64671;
    p25_add_65599 <= p25_add_65599_comb;
    p25_add_64308 <= p24_add_64308;
    p25_add_64552 <= p24_add_64552;
    p25_add_64290 <= p24_add_64290;
    p25_add_64289 <= p24_add_64289;
  end

  // ===== Pipe stage 26:
  wire [31:0] p26_add_65723_comb;
  wire [31:0] p26_and_65787_comb;
  wire [30:0] p26_add_65745_comb;
  wire [31:0] p26_add_65791_comb;
  wire [31:0] p26_add_65809_comb;
  wire [31:0] p26_add_65769_comb;
  wire [31:0] p26_add_65750_comb;
  wire [31:0] p26_add_65751_comb;
  wire [31:0] p26_add_65792_comb;
  wire [31:0] p26_add_65844_comb;
  wire [31:0] p26_add_65827_comb;
  wire [31:0] p26_add_65810_comb;
  wire [31:0] p26_add_65770_comb;
  wire [31:0] p26_add_65752_comb;
  assign p26_add_65723_comb = p25_add_65242 + p25_add_65599;
  assign p26_and_65787_comb = p25_add_65638 & p25_add_65519;
  assign p26_add_65745_comb = p25_add_64671[31:1] + 31'h3b7c_c46d;
  assign p26_add_65791_comb = {p25_add_65638[1:0] ^ p25_add_65638[12:11] ^ p25_add_65638[21:20], p25_add_65638[31:21] ^ p25_add_65638[10:0] ^ p25_add_65638[19:9], p25_add_65638[20:12] ^ p25_add_65638[31:23] ^ p25_add_65638[8:0], p25_add_65638[11:2] ^ p25_add_65638[22:13] ^ p25_add_65638[31:22]} + (p26_and_65787_comb ^ p25_add_65638 & p25_add_65342 ^ p25_and_65633);
  assign p26_add_65809_comb = p25_add_65616 + {p25_add_65029[16:7] ^ p25_add_65029[18:9], p25_add_65029[6:0] ^ p25_add_65029[8:2] ^ p25_add_65029[31:25], p25_add_65029[31:30] ^ p25_add_65029[1:0] ^ p25_add_65029[24:23], p25_add_65029[29:17] ^ p25_add_65029[31:19] ^ p25_add_65029[22:10]};
  assign p26_add_65769_comb = p25_add_64289 + {p25_add_65616[16:7] ^ p25_add_65616[18:9], p25_add_65616[6:0] ^ p25_add_65616[8:2] ^ p25_add_65616[31:25], p25_add_65616[31:30] ^ p25_add_65616[1:0] ^ p25_add_65616[24:23], p25_add_65616[29:17] ^ p25_add_65616[31:19] ^ p25_add_65616[22:10]};
  assign p26_add_65750_comb = {p26_add_65723_comb[5:0] ^ p26_add_65723_comb[10:5] ^ p26_add_65723_comb[24:19], p26_add_65723_comb[31:27] ^ p26_add_65723_comb[4:0] ^ p26_add_65723_comb[18:14], p26_add_65723_comb[26:13] ^ p26_add_65723_comb[31:18] ^ p26_add_65723_comb[13:0], p26_add_65723_comb[12:6] ^ p26_add_65723_comb[17:11] ^ p26_add_65723_comb[31:25]} + p25_add_65319;
  assign p26_add_65751_comb = (p26_add_65723_comb & p25_add_65570 ^ ~(p26_add_65723_comb | ~p25_add_65468)) + {p26_add_65745_comb, p25_add_64671[0]};
  assign p26_add_65792_comb = p25_add_65599 + p26_add_65791_comb;
  assign p26_add_65844_comb = {p25_add_64552[6:4] ^ p25_add_64552[17:15], p25_add_64552[3:0] ^ p25_add_64552[14:11] ^ p25_add_64552[31:28], p25_add_64552[31:21] ^ p25_add_64552[10:0] ^ p25_add_64552[27:17], p25_add_64552[20:7] ^ p25_add_64552[31:18] ^ p25_add_64552[16:3]} + p25_add_64290;
  assign p26_add_65827_comb = {p25_add_64290[6:4] ^ p25_add_64290[17:15], p25_add_64290[3:0] ^ p25_add_64290[14:11] ^ p25_add_64290[31:28], p25_add_64290[31:21] ^ p25_add_64290[10:0] ^ p25_add_64290[27:17], p25_add_64290[20:7] ^ p25_add_64290[31:18] ^ p25_add_64290[16:3]} + p25_add_64289;
  assign p26_add_65810_comb = p25_add_64325 + p26_add_65809_comb;
  assign p26_add_65770_comb = p25_add_64111 + p26_add_65769_comb;
  assign p26_add_65752_comb = p26_add_65750_comb + p26_add_65751_comb;

  // Registers for pipe stage 26:
  reg [31:0] p26_add_65468;
  reg [31:0] p26_add_65570;
  reg [31:0] p26_add_65723;
  reg [31:0] p26_add_65342;
  reg [31:0] p26_add_65519;
  reg [31:0] p26_add_65638;
  reg [31:0] p26_and_65787;
  reg [31:0] p26_add_65792;
  reg [31:0] p26_add_65844;
  reg [31:0] p26_add_65827;
  reg [31:0] p26_add_65672;
  reg [31:0] p26_add_65655;
  reg [31:0] p26_add_64810;
  reg [31:0] p26_add_65810;
  reg [31:0] p26_add_64179;
  reg [31:0] p26_add_65029;
  reg [31:0] p26_add_64145;
  reg [31:0] p26_add_64928;
  reg [31:0] p26_add_65770;
  reg [31:0] p26_add_64793;
  reg [31:0] p26_add_65616;
  reg [31:0] p26_add_65752;
  reg [31:0] p26_add_64671;
  reg [31:0] p26_add_64308;
  reg [31:0] p26_add_64552;
  always_ff @ (posedge clk) begin
    p26_add_65468 <= p25_add_65468;
    p26_add_65570 <= p25_add_65570;
    p26_add_65723 <= p26_add_65723_comb;
    p26_add_65342 <= p25_add_65342;
    p26_add_65519 <= p25_add_65519;
    p26_add_65638 <= p25_add_65638;
    p26_and_65787 <= p26_and_65787_comb;
    p26_add_65792 <= p26_add_65792_comb;
    p26_add_65844 <= p26_add_65844_comb;
    p26_add_65827 <= p26_add_65827_comb;
    p26_add_65672 <= p25_add_65672;
    p26_add_65655 <= p25_add_65655;
    p26_add_64810 <= p25_add_64810;
    p26_add_65810 <= p26_add_65810_comb;
    p26_add_64179 <= p25_add_64179;
    p26_add_65029 <= p25_add_65029;
    p26_add_64145 <= p25_add_64145;
    p26_add_64928 <= p25_add_64928;
    p26_add_65770 <= p26_add_65770_comb;
    p26_add_64793 <= p25_add_64793;
    p26_add_65616 <= p25_add_65616;
    p26_add_65752 <= p26_add_65752_comb;
    p26_add_64671 <= p25_add_64671;
    p26_add_64308 <= p25_add_64308;
    p26_add_64552 <= p25_add_64552;
  end

  // ===== Pipe stage 27:
  wire [31:0] p27_add_65895_comb;
  wire [31:0] p27_and_65942_comb;
  wire [30:0] p27_add_65917_comb;
  wire [31:0] p27_add_65946_comb;
  wire [31:0] p27_add_65982_comb;
  wire [31:0] p27_add_65964_comb;
  wire [31:0] p27_add_65922_comb;
  wire [31:0] p27_add_65923_comb;
  wire [31:0] p27_add_65925_comb;
  wire [31:0] p27_add_65947_comb;
  wire [31:0] p27_add_66017_comb;
  wire [31:0] p27_add_66000_comb;
  wire [31:0] p27_add_65983_comb;
  wire [31:0] p27_add_65965_comb;
  wire [31:0] p27_add_65924_comb;
  assign p27_add_65895_comb = p26_add_65342 + p26_add_65752;
  assign p27_and_65942_comb = p26_add_65792 & p26_add_65638;
  assign p27_add_65917_comb = p26_add_65616[31:1] + 31'h4c1f_28a9;
  assign p27_add_65946_comb = {p26_add_65792[1:0] ^ p26_add_65792[12:11] ^ p26_add_65792[21:20], p26_add_65792[31:21] ^ p26_add_65792[10:0] ^ p26_add_65792[19:9], p26_add_65792[20:12] ^ p26_add_65792[31:23] ^ p26_add_65792[8:0], p26_add_65792[11:2] ^ p26_add_65792[22:13] ^ p26_add_65792[31:22]} + (p27_and_65942_comb ^ p26_add_65792 & p26_add_65519 ^ p26_and_65787);
  assign p27_add_65982_comb = p26_add_65770 + {p26_add_65810[16:7] ^ p26_add_65810[18:9], p26_add_65810[6:0] ^ p26_add_65810[8:2] ^ p26_add_65810[31:25], p26_add_65810[31:30] ^ p26_add_65810[1:0] ^ p26_add_65810[24:23], p26_add_65810[29:17] ^ p26_add_65810[31:19] ^ p26_add_65810[22:10]};
  assign p27_add_65964_comb = p26_add_64552 + {p26_add_65770[16:7] ^ p26_add_65770[18:9], p26_add_65770[6:0] ^ p26_add_65770[8:2] ^ p26_add_65770[31:25], p26_add_65770[31:30] ^ p26_add_65770[1:0] ^ p26_add_65770[24:23], p26_add_65770[29:17] ^ p26_add_65770[31:19] ^ p26_add_65770[22:10]};
  assign p27_add_65922_comb = {p27_add_65895_comb[5:0] ^ p27_add_65895_comb[10:5] ^ p27_add_65895_comb[24:19], p27_add_65895_comb[31:27] ^ p27_add_65895_comb[4:0] ^ p27_add_65895_comb[18:14], p27_add_65895_comb[26:13] ^ p27_add_65895_comb[31:18] ^ p27_add_65895_comb[13:0], p27_add_65895_comb[12:6] ^ p27_add_65895_comb[17:11] ^ p27_add_65895_comb[31:25]} + p26_add_65468;
  assign p27_add_65923_comb = (p27_add_65895_comb & p26_add_65723 ^ ~(p27_add_65895_comb | ~p26_add_65570)) + {p27_add_65917_comb, p26_add_65616[0]};
  assign p27_add_65925_comb = p26_add_65570 + p26_add_64793;
  assign p27_add_65947_comb = p26_add_65752 + p27_add_65946_comb;
  assign p27_add_66017_comb = {p26_add_64671[6:4] ^ p26_add_64671[17:15], p26_add_64671[3:0] ^ p26_add_64671[14:11] ^ p26_add_64671[31:28], p26_add_64671[31:21] ^ p26_add_64671[10:0] ^ p26_add_64671[27:17], p26_add_64671[20:7] ^ p26_add_64671[31:18] ^ p26_add_64671[16:3]} + p26_add_64308;
  assign p27_add_66000_comb = {p26_add_64308[6:4] ^ p26_add_64308[17:15], p26_add_64308[3:0] ^ p26_add_64308[14:11] ^ p26_add_64308[31:28], p26_add_64308[31:21] ^ p26_add_64308[10:0] ^ p26_add_64308[27:17], p26_add_64308[20:7] ^ p26_add_64308[31:18] ^ p26_add_64308[16:3]} + p26_add_64552;
  assign p27_add_65983_comb = p26_add_65655 + p27_add_65982_comb;
  assign p27_add_65965_comb = p26_add_64145 + p27_add_65964_comb;
  assign p27_add_65924_comb = p27_add_65922_comb + p27_add_65923_comb;

  // Registers for pipe stage 27:
  reg [31:0] p27_add_65723;
  reg [31:0] p27_add_65895;
  reg [31:0] p27_add_65519;
  reg [31:0] p27_add_65925;
  reg [31:0] p27_add_65638;
  reg [31:0] p27_add_65792;
  reg [31:0] p27_and_65942;
  reg [31:0] p27_add_65947;
  reg [31:0] p27_add_66017;
  reg [31:0] p27_add_66000;
  reg [31:0] p27_add_65844;
  reg [31:0] p27_add_65827;
  reg [31:0] p27_add_65672;
  reg [31:0] p27_add_65983;
  reg [31:0] p27_add_64810;
  reg [31:0] p27_add_65810;
  reg [31:0] p27_add_64179;
  reg [31:0] p27_add_65029;
  reg [31:0] p27_add_65965;
  reg [31:0] p27_add_64928;
  reg [31:0] p27_add_65770;
  reg [31:0] p27_add_64793;
  reg [31:0] p27_add_65924;
  reg [31:0] p27_add_65616;
  reg [31:0] p27_add_64671;
  always_ff @ (posedge clk) begin
    p27_add_65723 <= p26_add_65723;
    p27_add_65895 <= p27_add_65895_comb;
    p27_add_65519 <= p26_add_65519;
    p27_add_65925 <= p27_add_65925_comb;
    p27_add_65638 <= p26_add_65638;
    p27_add_65792 <= p26_add_65792;
    p27_and_65942 <= p27_and_65942_comb;
    p27_add_65947 <= p27_add_65947_comb;
    p27_add_66017 <= p27_add_66017_comb;
    p27_add_66000 <= p27_add_66000_comb;
    p27_add_65844 <= p26_add_65844;
    p27_add_65827 <= p26_add_65827;
    p27_add_65672 <= p26_add_65672;
    p27_add_65983 <= p27_add_65983_comb;
    p27_add_64810 <= p26_add_64810;
    p27_add_65810 <= p26_add_65810;
    p27_add_64179 <= p26_add_64179;
    p27_add_65029 <= p26_add_65029;
    p27_add_65965 <= p27_add_65965_comb;
    p27_add_64928 <= p26_add_64928;
    p27_add_65770 <= p26_add_65770;
    p27_add_64793 <= p26_add_64793;
    p27_add_65924 <= p27_add_65924_comb;
    p27_add_65616 <= p26_add_65616;
    p27_add_64671 <= p26_add_64671;
  end

  // ===== Pipe stage 28:
  wire [31:0] p28_add_66068_comb;
  wire [31:0] p28_and_66109_comb;
  wire [31:0] p28_add_66113_comb;
  wire [31:0] p28_add_66090_comb;
  wire [31:0] p28_add_66149_comb;
  wire [31:0] p28_add_66131_comb;
  wire [31:0] p28_add_66114_comb;
  wire [31:0] p28_add_66092_comb;
  wire [31:0] p28_add_66184_comb;
  wire [31:0] p28_add_66167_comb;
  wire [31:0] p28_add_66150_comb;
  wire [31:0] p28_add_66132_comb;
  assign p28_add_66068_comb = p27_add_65519 + p27_add_65924;
  assign p28_and_66109_comb = p27_add_65947 & p27_add_65792;
  assign p28_add_66113_comb = {p27_add_65947[1:0] ^ p27_add_65947[12:11] ^ p27_add_65947[21:20], p27_add_65947[31:21] ^ p27_add_65947[10:0] ^ p27_add_65947[19:9], p27_add_65947[20:12] ^ p27_add_65947[31:23] ^ p27_add_65947[8:0], p27_add_65947[11:2] ^ p27_add_65947[22:13] ^ p27_add_65947[31:22]} + (p28_and_66109_comb ^ p27_add_65947 & p27_add_65638 ^ p27_and_65942);
  assign p28_add_66090_comb = {p28_add_66068_comb[5:0] ^ p28_add_66068_comb[10:5] ^ p28_add_66068_comb[24:19], p28_add_66068_comb[31:27] ^ p28_add_66068_comb[4:0] ^ p28_add_66068_comb[18:14], p28_add_66068_comb[26:13] ^ p28_add_66068_comb[31:18] ^ p28_add_66068_comb[13:0], p28_add_66068_comb[12:6] ^ p28_add_66068_comb[17:11] ^ p28_add_66068_comb[31:25]} + (p28_add_66068_comb & p27_add_65895 ^ ~(p28_add_66068_comb | ~p27_add_65723));
  assign p28_add_66149_comb = p27_add_65965 + {p27_add_65983[16:7] ^ p27_add_65983[18:9], p27_add_65983[6:0] ^ p27_add_65983[8:2] ^ p27_add_65983[31:25], p27_add_65983[31:30] ^ p27_add_65983[1:0] ^ p27_add_65983[24:23], p27_add_65983[29:17] ^ p27_add_65983[31:19] ^ p27_add_65983[22:10]};
  assign p28_add_66131_comb = p27_add_64671 + {p27_add_65965[16:7] ^ p27_add_65965[18:9], p27_add_65965[6:0] ^ p27_add_65965[8:2] ^ p27_add_65965[31:25], p27_add_65965[31:30] ^ p27_add_65965[1:0] ^ p27_add_65965[24:23], p27_add_65965[29:17] ^ p27_add_65965[31:19] ^ p27_add_65965[22:10]};
  assign p28_add_66114_comb = p27_add_65924 + p28_add_66113_comb;
  assign p28_add_66092_comb = p28_add_66090_comb + 32'ha831_c66d;
  assign p28_add_66184_comb = {p27_add_64793[6:4] ^ p27_add_64793[17:15], p27_add_64793[3:0] ^ p27_add_64793[14:11] ^ p27_add_64793[31:28], p27_add_64793[31:21] ^ p27_add_64793[10:0] ^ p27_add_64793[27:17], p27_add_64793[20:7] ^ p27_add_64793[31:18] ^ p27_add_64793[16:3]} + p27_add_65616;
  assign p28_add_66167_comb = {p27_add_65616[6:4] ^ p27_add_65616[17:15], p27_add_65616[3:0] ^ p27_add_65616[14:11] ^ p27_add_65616[31:28], p27_add_65616[31:21] ^ p27_add_65616[10:0] ^ p27_add_65616[27:17], p27_add_65616[20:7] ^ p27_add_65616[31:18] ^ p27_add_65616[16:3]} + p27_add_64671;
  assign p28_add_66150_comb = p27_add_65827 + p28_add_66149_comb;
  assign p28_add_66132_comb = p27_add_64179 + p28_add_66131_comb;

  // Registers for pipe stage 28:
  reg [31:0] p28_add_65723;
  reg [31:0] p28_add_65895;
  reg [31:0] p28_add_66068;
  reg [31:0] p28_add_65925;
  reg [31:0] p28_add_65638;
  reg [31:0] p28_add_65792;
  reg [31:0] p28_add_65947;
  reg [31:0] p28_and_66109;
  reg [31:0] p28_add_66114;
  reg [31:0] p28_add_66092;
  reg [31:0] p28_add_66184;
  reg [31:0] p28_add_66167;
  reg [31:0] p28_add_66017;
  reg [31:0] p28_add_66000;
  reg [31:0] p28_add_65844;
  reg [31:0] p28_add_66150;
  reg [31:0] p28_add_65672;
  reg [31:0] p28_add_65983;
  reg [31:0] p28_add_64810;
  reg [31:0] p28_add_65810;
  reg [31:0] p28_add_66132;
  reg [31:0] p28_add_65029;
  reg [31:0] p28_add_65965;
  reg [31:0] p28_add_64928;
  reg [31:0] p28_add_65770;
  reg [31:0] p28_add_64793;
  always_ff @ (posedge clk) begin
    p28_add_65723 <= p27_add_65723;
    p28_add_65895 <= p27_add_65895;
    p28_add_66068 <= p28_add_66068_comb;
    p28_add_65925 <= p27_add_65925;
    p28_add_65638 <= p27_add_65638;
    p28_add_65792 <= p27_add_65792;
    p28_add_65947 <= p27_add_65947;
    p28_and_66109 <= p28_and_66109_comb;
    p28_add_66114 <= p28_add_66114_comb;
    p28_add_66092 <= p28_add_66092_comb;
    p28_add_66184 <= p28_add_66184_comb;
    p28_add_66167 <= p28_add_66167_comb;
    p28_add_66017 <= p27_add_66017;
    p28_add_66000 <= p27_add_66000;
    p28_add_65844 <= p27_add_65844;
    p28_add_66150 <= p28_add_66150_comb;
    p28_add_65672 <= p27_add_65672;
    p28_add_65983 <= p27_add_65983;
    p28_add_64810 <= p27_add_64810;
    p28_add_65810 <= p27_add_65810;
    p28_add_66132 <= p28_add_66132_comb;
    p28_add_65029 <= p27_add_65029;
    p28_add_65965 <= p27_add_65965;
    p28_add_64928 <= p27_add_64928;
    p28_add_65770 <= p27_add_65770;
    p28_add_64793 <= p27_add_64793;
  end

  // ===== Pipe stage 29:
  wire [31:0] p29_add_66237_comb;
  wire [31:0] p29_add_66238_comb;
  wire [31:0] p29_and_66284_comb;
  wire [28:0] p29_add_66260_comb;
  wire [31:0] p29_add_66288_comb;
  wire [31:0] p29_add_66324_comb;
  wire [31:0] p29_add_66306_comb;
  wire [31:0] p29_add_66267_comb;
  wire [31:0] p29_add_66289_comb;
  wire [31:0] p29_add_66359_comb;
  wire [31:0] p29_add_66342_comb;
  wire [31:0] p29_add_66325_comb;
  wire [31:0] p29_add_66307_comb;
  wire [31:0] p29_add_66265_comb;
  wire [31:0] p29_add_66266_comb;
  assign p29_add_66237_comb = p28_add_66092 + p28_add_65925;
  assign p29_add_66238_comb = p28_add_65638 + p29_add_66237_comb;
  assign p29_and_66284_comb = p28_add_66114 & p28_add_65947;
  assign p29_add_66260_comb = p28_add_65770[31:3] + 29'h1600_64f9;
  assign p29_add_66288_comb = {p28_add_66114[1:0] ^ p28_add_66114[12:11] ^ p28_add_66114[21:20], p28_add_66114[31:21] ^ p28_add_66114[10:0] ^ p28_add_66114[19:9], p28_add_66114[20:12] ^ p28_add_66114[31:23] ^ p28_add_66114[8:0], p28_add_66114[11:2] ^ p28_add_66114[22:13] ^ p28_add_66114[31:22]} + (p29_and_66284_comb ^ p28_add_66114 & p28_add_65792 ^ p28_and_66109);
  assign p29_add_66324_comb = p28_add_66132 + {p28_add_66150[16:7] ^ p28_add_66150[18:9], p28_add_66150[6:0] ^ p28_add_66150[8:2] ^ p28_add_66150[31:25], p28_add_66150[31:30] ^ p28_add_66150[1:0] ^ p28_add_66150[24:23], p28_add_66150[29:17] ^ p28_add_66150[31:19] ^ p28_add_66150[22:10]};
  assign p29_add_66306_comb = p28_add_64793 + {p28_add_66132[16:7] ^ p28_add_66132[18:9], p28_add_66132[6:0] ^ p28_add_66132[8:2] ^ p28_add_66132[31:25], p28_add_66132[31:30] ^ p28_add_66132[1:0] ^ p28_add_66132[24:23], p28_add_66132[29:17] ^ p28_add_66132[31:19] ^ p28_add_66132[22:10]};
  assign p29_add_66267_comb = p28_add_65895 + p28_add_64928;
  assign p29_add_66289_comb = p29_add_66237_comb + p29_add_66288_comb;
  assign p29_add_66359_comb = {p28_add_64928[6:4] ^ p28_add_64928[17:15], p28_add_64928[3:0] ^ p28_add_64928[14:11] ^ p28_add_64928[31:28], p28_add_64928[31:21] ^ p28_add_64928[10:0] ^ p28_add_64928[27:17], p28_add_64928[20:7] ^ p28_add_64928[31:18] ^ p28_add_64928[16:3]} + p28_add_65770;
  assign p29_add_66342_comb = {p28_add_65770[6:4] ^ p28_add_65770[17:15], p28_add_65770[3:0] ^ p28_add_65770[14:11] ^ p28_add_65770[31:28], p28_add_65770[31:21] ^ p28_add_65770[10:0] ^ p28_add_65770[27:17], p28_add_65770[20:7] ^ p28_add_65770[31:18] ^ p28_add_65770[16:3]} + p28_add_64793;
  assign p29_add_66325_comb = p28_add_66000 + p29_add_66324_comb;
  assign p29_add_66307_comb = p28_add_64810 + p29_add_66306_comb;
  assign p29_add_66265_comb = {p29_add_66238_comb[5:0] ^ p29_add_66238_comb[10:5] ^ p29_add_66238_comb[24:19], p29_add_66238_comb[31:27] ^ p29_add_66238_comb[4:0] ^ p29_add_66238_comb[18:14], p29_add_66238_comb[26:13] ^ p29_add_66238_comb[31:18] ^ p29_add_66238_comb[13:0], p29_add_66238_comb[12:6] ^ p29_add_66238_comb[17:11] ^ p29_add_66238_comb[31:25]} + p28_add_65723;
  assign p29_add_66266_comb = (p29_add_66238_comb & p28_add_66068 ^ ~(p29_add_66238_comb | ~p28_add_65895)) + {p29_add_66260_comb, p28_add_65770[2:0]};

  // Registers for pipe stage 29:
  reg [31:0] p29_add_66068;
  reg [31:0] p29_add_66238;
  reg [31:0] p29_add_65792;
  reg [31:0] p29_add_66267;
  reg [31:0] p29_add_65947;
  reg [31:0] p29_add_66114;
  reg [31:0] p29_and_66284;
  reg [31:0] p29_add_66289;
  reg [31:0] p29_add_66359;
  reg [31:0] p29_add_66342;
  reg [31:0] p29_add_66184;
  reg [31:0] p29_add_66167;
  reg [31:0] p29_add_66017;
  reg [31:0] p29_add_66325;
  reg [31:0] p29_add_65844;
  reg [31:0] p29_add_66150;
  reg [31:0] p29_add_65672;
  reg [31:0] p29_add_65983;
  reg [31:0] p29_add_66307;
  reg [31:0] p29_add_65810;
  reg [31:0] p29_add_66132;
  reg [31:0] p29_add_65029;
  reg [31:0] p29_add_65965;
  reg [31:0] p29_add_64928;
  reg [31:0] p29_add_66265;
  reg [31:0] p29_add_66266;
  always_ff @ (posedge clk) begin
    p29_add_66068 <= p28_add_66068;
    p29_add_66238 <= p29_add_66238_comb;
    p29_add_65792 <= p28_add_65792;
    p29_add_66267 <= p29_add_66267_comb;
    p29_add_65947 <= p28_add_65947;
    p29_add_66114 <= p28_add_66114;
    p29_and_66284 <= p29_and_66284_comb;
    p29_add_66289 <= p29_add_66289_comb;
    p29_add_66359 <= p29_add_66359_comb;
    p29_add_66342 <= p29_add_66342_comb;
    p29_add_66184 <= p28_add_66184;
    p29_add_66167 <= p28_add_66167;
    p29_add_66017 <= p28_add_66017;
    p29_add_66325 <= p29_add_66325_comb;
    p29_add_65844 <= p28_add_65844;
    p29_add_66150 <= p28_add_66150;
    p29_add_65672 <= p28_add_65672;
    p29_add_65983 <= p28_add_65983;
    p29_add_66307 <= p29_add_66307_comb;
    p29_add_65810 <= p28_add_65810;
    p29_add_66132 <= p28_add_66132;
    p29_add_65029 <= p28_add_65029;
    p29_add_65965 <= p28_add_65965;
    p29_add_64928 <= p28_add_64928;
    p29_add_66265 <= p29_add_66265_comb;
    p29_add_66266 <= p29_add_66266_comb;
  end

  // ===== Pipe stage 30:
  wire [31:0] p30_add_66412_comb;
  wire [31:0] p30_add_66413_comb;
  wire [31:0] p30_and_66453_comb;
  wire [31:0] p30_add_66457_comb;
  wire [31:0] p30_add_66493_comb;
  wire [31:0] p30_add_66475_comb;
  wire [31:0] p30_add_66435_comb;
  wire [31:0] p30_add_66436_comb;
  wire [31:0] p30_add_66458_comb;
  wire [31:0] p30_add_66528_comb;
  wire [31:0] p30_add_66511_comb;
  wire [31:0] p30_add_66494_comb;
  wire [31:0] p30_add_66476_comb;
  assign p30_add_66412_comb = p29_add_66265 + p29_add_66266;
  assign p30_add_66413_comb = p29_add_65792 + p30_add_66412_comb;
  assign p30_and_66453_comb = p29_add_66289 & p29_add_66114;
  assign p30_add_66457_comb = {p29_add_66289[1:0] ^ p29_add_66289[12:11] ^ p29_add_66289[21:20], p29_add_66289[31:21] ^ p29_add_66289[10:0] ^ p29_add_66289[19:9], p29_add_66289[20:12] ^ p29_add_66289[31:23] ^ p29_add_66289[8:0], p29_add_66289[11:2] ^ p29_add_66289[22:13] ^ p29_add_66289[31:22]} + (p30_and_66453_comb ^ p29_add_66289 & p29_add_65947 ^ p29_and_66284);
  assign p30_add_66493_comb = p29_add_66307 + {p29_add_66325[16:7] ^ p29_add_66325[18:9], p29_add_66325[6:0] ^ p29_add_66325[8:2] ^ p29_add_66325[31:25], p29_add_66325[31:30] ^ p29_add_66325[1:0] ^ p29_add_66325[24:23], p29_add_66325[29:17] ^ p29_add_66325[31:19] ^ p29_add_66325[22:10]};
  assign p30_add_66475_comb = p29_add_64928 + {p29_add_66307[16:7] ^ p29_add_66307[18:9], p29_add_66307[6:0] ^ p29_add_66307[8:2] ^ p29_add_66307[31:25], p29_add_66307[31:30] ^ p29_add_66307[1:0] ^ p29_add_66307[24:23], p29_add_66307[29:17] ^ p29_add_66307[31:19] ^ p29_add_66307[22:10]};
  assign p30_add_66435_comb = {p30_add_66413_comb[5:0] ^ p30_add_66413_comb[10:5] ^ p30_add_66413_comb[24:19], p30_add_66413_comb[31:27] ^ p30_add_66413_comb[4:0] ^ p30_add_66413_comb[18:14], p30_add_66413_comb[26:13] ^ p30_add_66413_comb[31:18] ^ p30_add_66413_comb[13:0], p30_add_66413_comb[12:6] ^ p30_add_66413_comb[17:11] ^ p30_add_66413_comb[31:25]} + (p30_add_66413_comb & p29_add_66238 ^ ~(p30_add_66413_comb | ~p29_add_66068));
  assign p30_add_66436_comb = p29_add_66068 + p29_add_65965;
  assign p30_add_66458_comb = p30_add_66412_comb + p30_add_66457_comb;
  assign p30_add_66528_comb = {p29_add_65029[6:4] ^ p29_add_65029[17:15], p29_add_65029[3:0] ^ p29_add_65029[14:11] ^ p29_add_65029[31:28], p29_add_65029[31:21] ^ p29_add_65029[10:0] ^ p29_add_65029[27:17], p29_add_65029[20:7] ^ p29_add_65029[31:18] ^ p29_add_65029[16:3]} + p29_add_65965;
  assign p30_add_66511_comb = {p29_add_65965[6:4] ^ p29_add_65965[17:15], p29_add_65965[3:0] ^ p29_add_65965[14:11] ^ p29_add_65965[31:28], p29_add_65965[31:21] ^ p29_add_65965[10:0] ^ p29_add_65965[27:17], p29_add_65965[20:7] ^ p29_add_65965[31:18] ^ p29_add_65965[16:3]} + p29_add_64928;
  assign p30_add_66494_comb = p29_add_66167 + p30_add_66493_comb;
  assign p30_add_66476_comb = p29_add_65672 + p30_add_66475_comb;

  // Registers for pipe stage 30:
  reg [31:0] p30_add_66238;
  reg [31:0] p30_add_66413;
  reg [31:0] p30_add_66435;
  reg [31:0] p30_add_66267;
  reg [31:0] p30_add_65947;
  reg [31:0] p30_add_66436;
  reg [31:0] p30_add_66114;
  reg [31:0] p30_add_66289;
  reg [31:0] p30_and_66453;
  reg [31:0] p30_add_66458;
  reg [31:0] p30_add_66528;
  reg [31:0] p30_add_66511;
  reg [31:0] p30_add_66359;
  reg [31:0] p30_add_66342;
  reg [31:0] p30_add_66184;
  reg [31:0] p30_add_66494;
  reg [31:0] p30_add_66017;
  reg [31:0] p30_add_66325;
  reg [31:0] p30_add_65844;
  reg [31:0] p30_add_66150;
  reg [31:0] p30_add_66476;
  reg [31:0] p30_add_65983;
  reg [31:0] p30_add_66307;
  reg [31:0] p30_add_65810;
  reg [31:0] p30_add_66132;
  reg [31:0] p30_add_65029;
  always_ff @ (posedge clk) begin
    p30_add_66238 <= p29_add_66238;
    p30_add_66413 <= p30_add_66413_comb;
    p30_add_66435 <= p30_add_66435_comb;
    p30_add_66267 <= p29_add_66267;
    p30_add_65947 <= p29_add_65947;
    p30_add_66436 <= p30_add_66436_comb;
    p30_add_66114 <= p29_add_66114;
    p30_add_66289 <= p29_add_66289;
    p30_and_66453 <= p30_and_66453_comb;
    p30_add_66458 <= p30_add_66458_comb;
    p30_add_66528 <= p30_add_66528_comb;
    p30_add_66511 <= p30_add_66511_comb;
    p30_add_66359 <= p29_add_66359;
    p30_add_66342 <= p29_add_66342;
    p30_add_66184 <= p29_add_66184;
    p30_add_66494 <= p30_add_66494_comb;
    p30_add_66017 <= p29_add_66017;
    p30_add_66325 <= p29_add_66325;
    p30_add_65844 <= p29_add_65844;
    p30_add_66150 <= p29_add_66150;
    p30_add_66476 <= p30_add_66476_comb;
    p30_add_65983 <= p29_add_65983;
    p30_add_66307 <= p29_add_66307;
    p30_add_65810 <= p29_add_65810;
    p30_add_66132 <= p29_add_66132;
    p30_add_65029 <= p29_add_65029;
  end

  // ===== Pipe stage 31:
  wire [31:0] p31_and_66601_comb;
  wire [31:0] p31_add_66582_comb;
  wire [31:0] p31_add_66583_comb;
  wire [31:0] p31_add_66605_comb;
  wire [31:0] p31_add_66623_comb;
  wire [31:0] p31_add_66584_comb;
  wire [31:0] p31_add_66606_comb;
  wire [31:0] p31_add_66624_comb;
  assign p31_and_66601_comb = p30_add_66458 & p30_add_66289;
  assign p31_add_66582_comb = p30_add_66435 + 32'hbf59_7fc7;
  assign p31_add_66583_comb = p31_add_66582_comb + p30_add_66267;
  assign p31_add_66605_comb = {p30_add_66458[1:0] ^ p30_add_66458[12:11] ^ p30_add_66458[21:20], p30_add_66458[31:21] ^ p30_add_66458[10:0] ^ p30_add_66458[19:9], p30_add_66458[20:12] ^ p30_add_66458[31:23] ^ p30_add_66458[8:0], p30_add_66458[11:2] ^ p30_add_66458[22:13] ^ p30_add_66458[31:22]} + (p31_and_66601_comb ^ p30_add_66458 & p30_add_66114 ^ p30_and_66453);
  assign p31_add_66623_comb = p30_add_66476 + {p30_add_66494[16:7] ^ p30_add_66494[18:9], p30_add_66494[6:0] ^ p30_add_66494[8:2] ^ p30_add_66494[31:25], p30_add_66494[31:30] ^ p30_add_66494[1:0] ^ p30_add_66494[24:23], p30_add_66494[29:17] ^ p30_add_66494[31:19] ^ p30_add_66494[22:10]};
  assign p31_add_66584_comb = p30_add_65947 + p31_add_66583_comb;
  assign p31_add_66606_comb = p31_add_66583_comb + p31_add_66605_comb;
  assign p31_add_66624_comb = p30_add_66342 + p31_add_66623_comb;

  // Registers for pipe stage 31:
  reg [31:0] p31_add_66238;
  reg [31:0] p31_add_66413;
  reg [31:0] p31_add_66584;
  reg [31:0] p31_add_66436;
  reg [31:0] p31_add_66114;
  reg [31:0] p31_add_66289;
  reg [31:0] p31_add_66458;
  reg [31:0] p31_and_66601;
  reg [31:0] p31_add_66606;
  reg [31:0] p31_add_66528;
  reg [31:0] p31_add_66511;
  reg [31:0] p31_add_66359;
  reg [31:0] p31_add_66624;
  reg [31:0] p31_add_66184;
  reg [31:0] p31_add_66494;
  reg [31:0] p31_add_66017;
  reg [31:0] p31_add_66325;
  reg [31:0] p31_add_65844;
  reg [31:0] p31_add_66150;
  reg [31:0] p31_add_66476;
  reg [31:0] p31_add_65983;
  reg [31:0] p31_add_66307;
  reg [31:0] p31_add_65810;
  reg [31:0] p31_add_66132;
  reg [31:0] p31_add_65029;
  always_ff @ (posedge clk) begin
    p31_add_66238 <= p30_add_66238;
    p31_add_66413 <= p30_add_66413;
    p31_add_66584 <= p31_add_66584_comb;
    p31_add_66436 <= p30_add_66436;
    p31_add_66114 <= p30_add_66114;
    p31_add_66289 <= p30_add_66289;
    p31_add_66458 <= p30_add_66458;
    p31_and_66601 <= p31_and_66601_comb;
    p31_add_66606 <= p31_add_66606_comb;
    p31_add_66528 <= p30_add_66528;
    p31_add_66511 <= p30_add_66511;
    p31_add_66359 <= p30_add_66359;
    p31_add_66624 <= p31_add_66624_comb;
    p31_add_66184 <= p30_add_66184;
    p31_add_66494 <= p30_add_66494;
    p31_add_66017 <= p30_add_66017;
    p31_add_66325 <= p30_add_66325;
    p31_add_65844 <= p30_add_65844;
    p31_add_66150 <= p30_add_66150;
    p31_add_66476 <= p30_add_66476;
    p31_add_65983 <= p30_add_65983;
    p31_add_66307 <= p30_add_66307;
    p31_add_65810 <= p30_add_65810;
    p31_add_66132 <= p30_add_66132;
    p31_add_65029 <= p30_add_65029;
  end

  // ===== Pipe stage 32:
  wire [31:0] p32_add_66696_comb;
  wire [31:0] p32_add_66698_comb;
  wire [31:0] p32_add_66699_comb;
  wire [31:0] p32_add_66700_comb;
  assign p32_add_66696_comb = {p31_add_66584[5:0] ^ p31_add_66584[10:5] ^ p31_add_66584[24:19], p31_add_66584[31:27] ^ p31_add_66584[4:0] ^ p31_add_66584[18:14], p31_add_66584[26:13] ^ p31_add_66584[31:18] ^ p31_add_66584[13:0], p31_add_66584[12:6] ^ p31_add_66584[17:11] ^ p31_add_66584[31:25]} + (p31_add_66584 & p31_add_66413 ^ ~(p31_add_66584 | ~p31_add_66238));
  assign p32_add_66698_comb = p32_add_66696_comb + 32'hc6e0_0bf3;
  assign p32_add_66699_comb = p32_add_66698_comb + p31_add_66436;
  assign p32_add_66700_comb = p31_add_66238 + p31_add_65029;

  // Registers for pipe stage 32:
  reg [31:0] p32_add_66413;
  reg [31:0] p32_add_66584;
  reg [31:0] p32_add_66114;
  reg [31:0] p32_add_66699;
  reg [31:0] p32_add_66700;
  reg [31:0] p32_add_66289;
  reg [31:0] p32_add_66458;
  reg [31:0] p32_and_66601;
  reg [31:0] p32_add_66606;
  reg [31:0] p32_add_66528;
  reg [31:0] p32_add_66511;
  reg [31:0] p32_add_66359;
  reg [31:0] p32_add_66624;
  reg [31:0] p32_add_66184;
  reg [31:0] p32_add_66494;
  reg [31:0] p32_add_66017;
  reg [31:0] p32_add_66325;
  reg [31:0] p32_add_65844;
  reg [31:0] p32_add_66150;
  reg [31:0] p32_add_66476;
  reg [31:0] p32_add_65983;
  reg [31:0] p32_add_66307;
  reg [31:0] p32_add_65810;
  reg [31:0] p32_add_66132;
  reg [31:0] p32_add_65029;
  always_ff @ (posedge clk) begin
    p32_add_66413 <= p31_add_66413;
    p32_add_66584 <= p31_add_66584;
    p32_add_66114 <= p31_add_66114;
    p32_add_66699 <= p32_add_66699_comb;
    p32_add_66700 <= p32_add_66700_comb;
    p32_add_66289 <= p31_add_66289;
    p32_add_66458 <= p31_add_66458;
    p32_and_66601 <= p31_and_66601;
    p32_add_66606 <= p31_add_66606;
    p32_add_66528 <= p31_add_66528;
    p32_add_66511 <= p31_add_66511;
    p32_add_66359 <= p31_add_66359;
    p32_add_66624 <= p31_add_66624;
    p32_add_66184 <= p31_add_66184;
    p32_add_66494 <= p31_add_66494;
    p32_add_66017 <= p31_add_66017;
    p32_add_66325 <= p31_add_66325;
    p32_add_65844 <= p31_add_65844;
    p32_add_66150 <= p31_add_66150;
    p32_add_66476 <= p31_add_66476;
    p32_add_65983 <= p31_add_65983;
    p32_add_66307 <= p31_add_66307;
    p32_add_65810 <= p31_add_65810;
    p32_add_66132 <= p31_add_66132;
    p32_add_65029 <= p31_add_65029;
  end

  // ===== Pipe stage 33:
  wire [31:0] p33_add_66751_comb;
  wire [31:0] p33_and_66793_comb;
  wire [31:0] p33_add_66797_comb;
  wire [31:0] p33_add_66773_comb;
  wire [31:0] p33_add_66776_comb;
  wire [31:0] p33_add_66798_comb;
  wire [31:0] p33_add_66775_comb;
  assign p33_add_66751_comb = p32_add_66114 + p32_add_66699;
  assign p33_and_66793_comb = p32_add_66606 & p32_add_66458;
  assign p33_add_66797_comb = {p32_add_66606[1:0] ^ p32_add_66606[12:11] ^ p32_add_66606[21:20], p32_add_66606[31:21] ^ p32_add_66606[10:0] ^ p32_add_66606[19:9], p32_add_66606[20:12] ^ p32_add_66606[31:23] ^ p32_add_66606[8:0], p32_add_66606[11:2] ^ p32_add_66606[22:13] ^ p32_add_66606[31:22]} + (p33_and_66793_comb ^ p32_add_66606 & p32_add_66289 ^ p32_and_66601);
  assign p33_add_66773_comb = {p33_add_66751_comb[5:0] ^ p33_add_66751_comb[10:5] ^ p33_add_66751_comb[24:19], p33_add_66751_comb[31:27] ^ p33_add_66751_comb[4:0] ^ p33_add_66751_comb[18:14], p33_add_66751_comb[26:13] ^ p33_add_66751_comb[31:18] ^ p33_add_66751_comb[13:0], p33_add_66751_comb[12:6] ^ p33_add_66751_comb[17:11] ^ p33_add_66751_comb[31:25]} + (p33_add_66751_comb & p32_add_66584 ^ ~(p33_add_66751_comb | ~p32_add_66413));
  assign p33_add_66776_comb = p32_add_66413 + p32_add_66132;
  assign p33_add_66798_comb = p32_add_66699 + p33_add_66797_comb;
  assign p33_add_66775_comb = p33_add_66773_comb + 32'hd5a7_9147;

  // Registers for pipe stage 33:
  reg [31:0] p33_add_66584;
  reg [31:0] p33_add_66751;
  reg [31:0] p33_add_66700;
  reg [31:0] p33_add_66289;
  reg [31:0] p33_add_66776;
  reg [31:0] p33_add_66458;
  reg [31:0] p33_add_66606;
  reg [31:0] p33_and_66793;
  reg [31:0] p33_add_66798;
  reg [31:0] p33_add_66775;
  reg [31:0] p33_add_66528;
  reg [31:0] p33_add_66511;
  reg [31:0] p33_add_66359;
  reg [31:0] p33_add_66624;
  reg [31:0] p33_add_66184;
  reg [31:0] p33_add_66494;
  reg [31:0] p33_add_66017;
  reg [31:0] p33_add_66325;
  reg [31:0] p33_add_65844;
  reg [31:0] p33_add_66150;
  reg [31:0] p33_add_66476;
  reg [31:0] p33_add_65983;
  reg [31:0] p33_add_66307;
  reg [31:0] p33_add_65810;
  reg [31:0] p33_add_66132;
  reg [31:0] p33_add_65029;
  always_ff @ (posedge clk) begin
    p33_add_66584 <= p32_add_66584;
    p33_add_66751 <= p33_add_66751_comb;
    p33_add_66700 <= p32_add_66700;
    p33_add_66289 <= p32_add_66289;
    p33_add_66776 <= p33_add_66776_comb;
    p33_add_66458 <= p32_add_66458;
    p33_add_66606 <= p32_add_66606;
    p33_and_66793 <= p33_and_66793_comb;
    p33_add_66798 <= p33_add_66798_comb;
    p33_add_66775 <= p33_add_66775_comb;
    p33_add_66528 <= p32_add_66528;
    p33_add_66511 <= p32_add_66511;
    p33_add_66359 <= p32_add_66359;
    p33_add_66624 <= p32_add_66624;
    p33_add_66184 <= p32_add_66184;
    p33_add_66494 <= p32_add_66494;
    p33_add_66017 <= p32_add_66017;
    p33_add_66325 <= p32_add_66325;
    p33_add_65844 <= p32_add_65844;
    p33_add_66150 <= p32_add_66150;
    p33_add_66476 <= p32_add_66476;
    p33_add_65983 <= p32_add_65983;
    p33_add_66307 <= p32_add_66307;
    p33_add_65810 <= p32_add_65810;
    p33_add_66132 <= p32_add_66132;
    p33_add_65029 <= p32_add_65029;
  end

  // ===== Pipe stage 34:
  wire [31:0] p34_add_66851_comb;
  wire [31:0] p34_add_66852_comb;
  wire [31:0] p34_and_66892_comb;
  wire [31:0] p34_add_66896_comb;
  wire [31:0] p34_add_66874_comb;
  wire [31:0] p34_add_66875_comb;
  wire [31:0] p34_add_66897_comb;
  assign p34_add_66851_comb = p33_add_66775 + p33_add_66700;
  assign p34_add_66852_comb = p33_add_66289 + p34_add_66851_comb;
  assign p34_and_66892_comb = p33_add_66798 & p33_add_66606;
  assign p34_add_66896_comb = {p33_add_66798[1:0] ^ p33_add_66798[12:11] ^ p33_add_66798[21:20], p33_add_66798[31:21] ^ p33_add_66798[10:0] ^ p33_add_66798[19:9], p33_add_66798[20:12] ^ p33_add_66798[31:23] ^ p33_add_66798[8:0], p33_add_66798[11:2] ^ p33_add_66798[22:13] ^ p33_add_66798[31:22]} + (p34_and_66892_comb ^ p33_add_66798 & p33_add_66458 ^ p33_and_66793);
  assign p34_add_66874_comb = {p34_add_66852_comb[5:0] ^ p34_add_66852_comb[10:5] ^ p34_add_66852_comb[24:19], p34_add_66852_comb[31:27] ^ p34_add_66852_comb[4:0] ^ p34_add_66852_comb[18:14], p34_add_66852_comb[26:13] ^ p34_add_66852_comb[31:18] ^ p34_add_66852_comb[13:0], p34_add_66852_comb[12:6] ^ p34_add_66852_comb[17:11] ^ p34_add_66852_comb[31:25]} + (p34_add_66852_comb & p33_add_66751 ^ ~(p34_add_66852_comb | ~p33_add_66584));
  assign p34_add_66875_comb = p33_add_66584 + p33_add_65810;
  assign p34_add_66897_comb = p34_add_66851_comb + p34_add_66896_comb;

  // Registers for pipe stage 34:
  reg [31:0] p34_add_66751;
  reg [31:0] p34_add_66852;
  reg [31:0] p34_add_66874;
  reg [31:0] p34_add_66776;
  reg [31:0] p34_add_66458;
  reg [31:0] p34_add_66875;
  reg [31:0] p34_add_66606;
  reg [31:0] p34_add_66798;
  reg [31:0] p34_and_66892;
  reg [31:0] p34_add_66897;
  reg [31:0] p34_add_66528;
  reg [31:0] p34_add_66511;
  reg [31:0] p34_add_66359;
  reg [31:0] p34_add_66624;
  reg [31:0] p34_add_66184;
  reg [31:0] p34_add_66494;
  reg [31:0] p34_add_66017;
  reg [31:0] p34_add_66325;
  reg [31:0] p34_add_65844;
  reg [31:0] p34_add_66150;
  reg [31:0] p34_add_66476;
  reg [31:0] p34_add_65983;
  reg [31:0] p34_add_66307;
  reg [31:0] p34_add_65810;
  reg [31:0] p34_add_66132;
  reg [31:0] p34_add_65029;
  always_ff @ (posedge clk) begin
    p34_add_66751 <= p33_add_66751;
    p34_add_66852 <= p34_add_66852_comb;
    p34_add_66874 <= p34_add_66874_comb;
    p34_add_66776 <= p33_add_66776;
    p34_add_66458 <= p33_add_66458;
    p34_add_66875 <= p34_add_66875_comb;
    p34_add_66606 <= p33_add_66606;
    p34_add_66798 <= p33_add_66798;
    p34_and_66892 <= p34_and_66892_comb;
    p34_add_66897 <= p34_add_66897_comb;
    p34_add_66528 <= p33_add_66528;
    p34_add_66511 <= p33_add_66511;
    p34_add_66359 <= p33_add_66359;
    p34_add_66624 <= p33_add_66624;
    p34_add_66184 <= p33_add_66184;
    p34_add_66494 <= p33_add_66494;
    p34_add_66017 <= p33_add_66017;
    p34_add_66325 <= p33_add_66325;
    p34_add_65844 <= p33_add_65844;
    p34_add_66150 <= p33_add_66150;
    p34_add_66476 <= p33_add_66476;
    p34_add_65983 <= p33_add_65983;
    p34_add_66307 <= p33_add_66307;
    p34_add_65810 <= p33_add_65810;
    p34_add_66132 <= p33_add_66132;
    p34_add_65029 <= p33_add_65029;
  end

  // ===== Pipe stage 35:
  wire [31:0] p35_and_66970_comb;
  wire [31:0] p35_add_66951_comb;
  wire [31:0] p35_add_66952_comb;
  wire [31:0] p35_add_66974_comb;
  wire [31:0] p35_add_66953_comb;
  wire [31:0] p35_add_66975_comb;
  assign p35_and_66970_comb = p34_add_66897 & p34_add_66798;
  assign p35_add_66951_comb = p34_add_66874 + 32'h06ca_6351;
  assign p35_add_66952_comb = p35_add_66951_comb + p34_add_66776;
  assign p35_add_66974_comb = {p34_add_66897[1:0] ^ p34_add_66897[12:11] ^ p34_add_66897[21:20], p34_add_66897[31:21] ^ p34_add_66897[10:0] ^ p34_add_66897[19:9], p34_add_66897[20:12] ^ p34_add_66897[31:23] ^ p34_add_66897[8:0], p34_add_66897[11:2] ^ p34_add_66897[22:13] ^ p34_add_66897[31:22]} + (p35_and_66970_comb ^ p34_add_66897 & p34_add_66606 ^ p34_and_66892);
  assign p35_add_66953_comb = p34_add_66458 + p35_add_66952_comb;
  assign p35_add_66975_comb = p35_add_66952_comb + p35_add_66974_comb;

  // Registers for pipe stage 35:
  reg [31:0] p35_add_66751;
  reg [31:0] p35_add_66852;
  reg [31:0] p35_add_66953;
  reg [31:0] p35_add_66875;
  reg [31:0] p35_add_66606;
  reg [31:0] p35_add_66798;
  reg [31:0] p35_add_66897;
  reg [31:0] p35_and_66970;
  reg [31:0] p35_add_66975;
  reg [31:0] p35_add_66528;
  reg [31:0] p35_add_66511;
  reg [31:0] p35_add_66359;
  reg [31:0] p35_add_66624;
  reg [31:0] p35_add_66184;
  reg [31:0] p35_add_66494;
  reg [31:0] p35_add_66017;
  reg [31:0] p35_add_66325;
  reg [31:0] p35_add_65844;
  reg [31:0] p35_add_66150;
  reg [31:0] p35_add_66476;
  reg [31:0] p35_add_65983;
  reg [31:0] p35_add_66307;
  reg [31:0] p35_add_65810;
  reg [31:0] p35_add_66132;
  reg [31:0] p35_add_65029;
  always_ff @ (posedge clk) begin
    p35_add_66751 <= p34_add_66751;
    p35_add_66852 <= p34_add_66852;
    p35_add_66953 <= p35_add_66953_comb;
    p35_add_66875 <= p34_add_66875;
    p35_add_66606 <= p34_add_66606;
    p35_add_66798 <= p34_add_66798;
    p35_add_66897 <= p34_add_66897;
    p35_and_66970 <= p35_and_66970_comb;
    p35_add_66975 <= p35_add_66975_comb;
    p35_add_66528 <= p34_add_66528;
    p35_add_66511 <= p34_add_66511;
    p35_add_66359 <= p34_add_66359;
    p35_add_66624 <= p34_add_66624;
    p35_add_66184 <= p34_add_66184;
    p35_add_66494 <= p34_add_66494;
    p35_add_66017 <= p34_add_66017;
    p35_add_66325 <= p34_add_66325;
    p35_add_65844 <= p34_add_65844;
    p35_add_66150 <= p34_add_66150;
    p35_add_66476 <= p34_add_66476;
    p35_add_65983 <= p34_add_65983;
    p35_add_66307 <= p34_add_66307;
    p35_add_65810 <= p34_add_65810;
    p35_add_66132 <= p34_add_66132;
    p35_add_65029 <= p34_add_65029;
  end

  // ===== Pipe stage 36:
  wire [31:0] p36_add_67047_comb;
  wire [31:0] p36_add_67049_comb;
  wire [31:0] p36_add_67050_comb;
  wire [31:0] p36_add_67051_comb;
  assign p36_add_67047_comb = {p35_add_66953[5:0] ^ p35_add_66953[10:5] ^ p35_add_66953[24:19], p35_add_66953[31:27] ^ p35_add_66953[4:0] ^ p35_add_66953[18:14], p35_add_66953[26:13] ^ p35_add_66953[31:18] ^ p35_add_66953[13:0], p35_add_66953[12:6] ^ p35_add_66953[17:11] ^ p35_add_66953[31:25]} + (p35_add_66953 & p35_add_66852 ^ ~(p35_add_66953 | ~p35_add_66751));
  assign p36_add_67049_comb = p36_add_67047_comb + 32'h1429_2967;
  assign p36_add_67050_comb = p36_add_67049_comb + p35_add_66875;
  assign p36_add_67051_comb = p35_add_66751 + p35_add_66307;

  // Registers for pipe stage 36:
  reg [31:0] p36_add_66852;
  reg [31:0] p36_add_66953;
  reg [31:0] p36_add_66606;
  reg [31:0] p36_add_67050;
  reg [31:0] p36_add_67051;
  reg [31:0] p36_add_66798;
  reg [31:0] p36_add_66897;
  reg [31:0] p36_and_66970;
  reg [31:0] p36_add_66975;
  reg [31:0] p36_add_66528;
  reg [31:0] p36_add_66511;
  reg [31:0] p36_add_66359;
  reg [31:0] p36_add_66624;
  reg [31:0] p36_add_66184;
  reg [31:0] p36_add_66494;
  reg [31:0] p36_add_66017;
  reg [31:0] p36_add_66325;
  reg [31:0] p36_add_65844;
  reg [31:0] p36_add_66150;
  reg [31:0] p36_add_66476;
  reg [31:0] p36_add_65983;
  reg [31:0] p36_add_66307;
  reg [31:0] p36_add_65810;
  reg [31:0] p36_add_66132;
  reg [31:0] p36_add_65029;
  always_ff @ (posedge clk) begin
    p36_add_66852 <= p35_add_66852;
    p36_add_66953 <= p35_add_66953;
    p36_add_66606 <= p35_add_66606;
    p36_add_67050 <= p36_add_67050_comb;
    p36_add_67051 <= p36_add_67051_comb;
    p36_add_66798 <= p35_add_66798;
    p36_add_66897 <= p35_add_66897;
    p36_and_66970 <= p35_and_66970;
    p36_add_66975 <= p35_add_66975;
    p36_add_66528 <= p35_add_66528;
    p36_add_66511 <= p35_add_66511;
    p36_add_66359 <= p35_add_66359;
    p36_add_66624 <= p35_add_66624;
    p36_add_66184 <= p35_add_66184;
    p36_add_66494 <= p35_add_66494;
    p36_add_66017 <= p35_add_66017;
    p36_add_66325 <= p35_add_66325;
    p36_add_65844 <= p35_add_65844;
    p36_add_66150 <= p35_add_66150;
    p36_add_66476 <= p35_add_66476;
    p36_add_65983 <= p35_add_65983;
    p36_add_66307 <= p35_add_66307;
    p36_add_65810 <= p35_add_65810;
    p36_add_66132 <= p35_add_66132;
    p36_add_65029 <= p35_add_65029;
  end

  // ===== Pipe stage 37:
  wire [31:0] p37_add_67102_comb;
  wire [31:0] p37_and_67143_comb;
  wire [31:0] p37_add_67147_comb;
  wire [31:0] p37_add_67124_comb;
  wire [31:0] p37_add_67148_comb;
  wire [31:0] p37_add_67126_comb;
  assign p37_add_67102_comb = p36_add_66606 + p36_add_67050;
  assign p37_and_67143_comb = p36_add_66975 & p36_add_66897;
  assign p37_add_67147_comb = {p36_add_66975[1:0] ^ p36_add_66975[12:11] ^ p36_add_66975[21:20], p36_add_66975[31:21] ^ p36_add_66975[10:0] ^ p36_add_66975[19:9], p36_add_66975[20:12] ^ p36_add_66975[31:23] ^ p36_add_66975[8:0], p36_add_66975[11:2] ^ p36_add_66975[22:13] ^ p36_add_66975[31:22]} + (p37_and_67143_comb ^ p36_add_66975 & p36_add_66798 ^ p36_and_66970);
  assign p37_add_67124_comb = {p37_add_67102_comb[5:0] ^ p37_add_67102_comb[10:5] ^ p37_add_67102_comb[24:19], p37_add_67102_comb[31:27] ^ p37_add_67102_comb[4:0] ^ p37_add_67102_comb[18:14], p37_add_67102_comb[26:13] ^ p37_add_67102_comb[31:18] ^ p37_add_67102_comb[13:0], p37_add_67102_comb[12:6] ^ p37_add_67102_comb[17:11] ^ p37_add_67102_comb[31:25]} + (p37_add_67102_comb & p36_add_66953 ^ ~(p37_add_67102_comb | ~p36_add_66852));
  assign p37_add_67148_comb = p36_add_67050 + p37_add_67147_comb;
  assign p37_add_67126_comb = p37_add_67124_comb + 32'h27b7_0a85;

  // Registers for pipe stage 37:
  reg [31:0] p37_add_66852;
  reg [31:0] p37_add_66953;
  reg [31:0] p37_add_67102;
  reg [31:0] p37_add_67051;
  reg [31:0] p37_add_66798;
  reg [31:0] p37_add_66897;
  reg [31:0] p37_add_66975;
  reg [31:0] p37_and_67143;
  reg [31:0] p37_add_67148;
  reg [31:0] p37_add_67126;
  reg [31:0] p37_add_66528;
  reg [31:0] p37_add_66511;
  reg [31:0] p37_add_66359;
  reg [31:0] p37_add_66624;
  reg [31:0] p37_add_66184;
  reg [31:0] p37_add_66494;
  reg [31:0] p37_add_66017;
  reg [31:0] p37_add_66325;
  reg [31:0] p37_add_65844;
  reg [31:0] p37_add_66150;
  reg [31:0] p37_add_66476;
  reg [31:0] p37_add_65983;
  reg [31:0] p37_add_66307;
  reg [31:0] p37_add_65810;
  reg [31:0] p37_add_66132;
  reg [31:0] p37_add_65029;
  always_ff @ (posedge clk) begin
    p37_add_66852 <= p36_add_66852;
    p37_add_66953 <= p36_add_66953;
    p37_add_67102 <= p37_add_67102_comb;
    p37_add_67051 <= p36_add_67051;
    p37_add_66798 <= p36_add_66798;
    p37_add_66897 <= p36_add_66897;
    p37_add_66975 <= p36_add_66975;
    p37_and_67143 <= p37_and_67143_comb;
    p37_add_67148 <= p37_add_67148_comb;
    p37_add_67126 <= p37_add_67126_comb;
    p37_add_66528 <= p36_add_66528;
    p37_add_66511 <= p36_add_66511;
    p37_add_66359 <= p36_add_66359;
    p37_add_66624 <= p36_add_66624;
    p37_add_66184 <= p36_add_66184;
    p37_add_66494 <= p36_add_66494;
    p37_add_66017 <= p36_add_66017;
    p37_add_66325 <= p36_add_66325;
    p37_add_65844 <= p36_add_65844;
    p37_add_66150 <= p36_add_66150;
    p37_add_66476 <= p36_add_66476;
    p37_add_65983 <= p36_add_65983;
    p37_add_66307 <= p36_add_66307;
    p37_add_65810 <= p36_add_65810;
    p37_add_66132 <= p36_add_66132;
    p37_add_65029 <= p36_add_65029;
  end

  // ===== Pipe stage 38:
  wire [31:0] p38_add_67201_comb;
  wire [31:0] p38_add_67202_comb;
  wire [31:0] p38_and_67247_comb;
  wire [28:0] p38_add_67224_comb;
  wire [31:0] p38_add_67251_comb;
  wire [31:0] p38_add_67252_comb;
  wire [31:0] p38_add_67229_comb;
  wire [31:0] p38_add_67230_comb;
  assign p38_add_67201_comb = p37_add_67126 + p37_add_67051;
  assign p38_add_67202_comb = p37_add_66798 + p38_add_67201_comb;
  assign p38_and_67247_comb = p37_add_67148 & p37_add_66975;
  assign p38_add_67224_comb = p37_add_65983[31:3] + 29'h05c3_6427;
  assign p38_add_67251_comb = {p37_add_67148[1:0] ^ p37_add_67148[12:11] ^ p37_add_67148[21:20], p37_add_67148[31:21] ^ p37_add_67148[10:0] ^ p37_add_67148[19:9], p37_add_67148[20:12] ^ p37_add_67148[31:23] ^ p37_add_67148[8:0], p37_add_67148[11:2] ^ p37_add_67148[22:13] ^ p37_add_67148[31:22]} + (p38_and_67247_comb ^ p37_add_67148 & p37_add_66897 ^ p37_and_67143);
  assign p38_add_67252_comb = p38_add_67201_comb + p38_add_67251_comb;
  assign p38_add_67229_comb = {p38_add_67202_comb[5:0] ^ p38_add_67202_comb[10:5] ^ p38_add_67202_comb[24:19], p38_add_67202_comb[31:27] ^ p38_add_67202_comb[4:0] ^ p38_add_67202_comb[18:14], p38_add_67202_comb[26:13] ^ p38_add_67202_comb[31:18] ^ p38_add_67202_comb[13:0], p38_add_67202_comb[12:6] ^ p38_add_67202_comb[17:11] ^ p38_add_67202_comb[31:25]} + p37_add_66852;
  assign p38_add_67230_comb = (p38_add_67202_comb & p37_add_67102 ^ ~(p38_add_67202_comb | ~p37_add_66953)) + {p38_add_67224_comb, p37_add_65983[2:0]};

  // Registers for pipe stage 38:
  reg [31:0] p38_add_66953;
  reg [31:0] p38_add_67102;
  reg [31:0] p38_add_67202;
  reg [31:0] p38_add_66897;
  reg [31:0] p38_add_66975;
  reg [31:0] p38_add_67148;
  reg [31:0] p38_and_67247;
  reg [31:0] p38_add_67252;
  reg [31:0] p38_add_66528;
  reg [31:0] p38_add_66511;
  reg [31:0] p38_add_66359;
  reg [31:0] p38_add_66624;
  reg [31:0] p38_add_66184;
  reg [31:0] p38_add_66494;
  reg [31:0] p38_add_66017;
  reg [31:0] p38_add_66325;
  reg [31:0] p38_add_65844;
  reg [31:0] p38_add_66150;
  reg [31:0] p38_add_66476;
  reg [31:0] p38_add_67229;
  reg [31:0] p38_add_67230;
  reg [31:0] p38_add_65983;
  reg [31:0] p38_add_66307;
  reg [31:0] p38_add_65810;
  reg [31:0] p38_add_66132;
  reg [31:0] p38_add_65029;
  always_ff @ (posedge clk) begin
    p38_add_66953 <= p37_add_66953;
    p38_add_67102 <= p37_add_67102;
    p38_add_67202 <= p38_add_67202_comb;
    p38_add_66897 <= p37_add_66897;
    p38_add_66975 <= p37_add_66975;
    p38_add_67148 <= p37_add_67148;
    p38_and_67247 <= p38_and_67247_comb;
    p38_add_67252 <= p38_add_67252_comb;
    p38_add_66528 <= p37_add_66528;
    p38_add_66511 <= p37_add_66511;
    p38_add_66359 <= p37_add_66359;
    p38_add_66624 <= p37_add_66624;
    p38_add_66184 <= p37_add_66184;
    p38_add_66494 <= p37_add_66494;
    p38_add_66017 <= p37_add_66017;
    p38_add_66325 <= p37_add_66325;
    p38_add_65844 <= p37_add_65844;
    p38_add_66150 <= p37_add_66150;
    p38_add_66476 <= p37_add_66476;
    p38_add_67229 <= p38_add_67229_comb;
    p38_add_67230 <= p38_add_67230_comb;
    p38_add_65983 <= p37_add_65983;
    p38_add_66307 <= p37_add_66307;
    p38_add_65810 <= p37_add_65810;
    p38_add_66132 <= p37_add_66132;
    p38_add_65029 <= p37_add_65029;
  end

  // ===== Pipe stage 39:
  wire [31:0] p39_add_67305_comb;
  wire [31:0] p39_add_67306_comb;
  wire [31:0] p39_and_67369_comb;
  wire [29:0] p39_add_67328_comb;
  wire [31:0] p39_add_67373_comb;
  wire [31:0] p39_add_67351_comb;
  wire [31:0] p39_add_67349_comb;
  wire [31:0] p39_add_67374_comb;
  wire [31:0] p39_add_67408_comb;
  wire [31:0] p39_add_67391_comb;
  wire [31:0] p39_add_67352_comb;
  wire [31:0] p39_add_67333_comb;
  wire [31:0] p39_add_67334_comb;
  assign p39_add_67305_comb = p38_add_67229 + p38_add_67230;
  assign p39_add_67306_comb = p38_add_66897 + p39_add_67305_comb;
  assign p39_and_67369_comb = p38_add_67252 & p38_add_67148;
  assign p39_add_67328_comb = p38_add_66476[31:2] + 30'h134b_1b7f;
  assign p39_add_67373_comb = {p38_add_67252[1:0] ^ p38_add_67252[12:11] ^ p38_add_67252[21:20], p38_add_67252[31:21] ^ p38_add_67252[10:0] ^ p38_add_67252[19:9], p38_add_67252[20:12] ^ p38_add_67252[31:23] ^ p38_add_67252[8:0], p38_add_67252[11:2] ^ p38_add_67252[22:13] ^ p38_add_67252[31:22]} + (p39_and_67369_comb ^ p38_add_67252 & p38_add_66975 ^ p38_and_67247);
  assign p39_add_67351_comb = p38_add_65029 + {p38_add_66476[16:7] ^ p38_add_66476[18:9], p38_add_66476[6:0] ^ p38_add_66476[8:2] ^ p38_add_66476[31:25], p38_add_66476[31:30] ^ p38_add_66476[1:0] ^ p38_add_66476[24:23], p38_add_66476[29:17] ^ p38_add_66476[31:19] ^ p38_add_66476[22:10]};
  assign p39_add_67349_comb = p38_add_67102 + p38_add_66150;
  assign p39_add_67374_comb = p39_add_67305_comb + p39_add_67373_comb;
  assign p39_add_67408_comb = {p38_add_65810[6:4] ^ p38_add_65810[17:15], p38_add_65810[3:0] ^ p38_add_65810[14:11] ^ p38_add_65810[31:28], p38_add_65810[31:21] ^ p38_add_65810[10:0] ^ p38_add_65810[27:17], p38_add_65810[20:7] ^ p38_add_65810[31:18] ^ p38_add_65810[16:3]} + p38_add_66132;
  assign p39_add_67391_comb = {p38_add_66132[6:4] ^ p38_add_66132[17:15], p38_add_66132[3:0] ^ p38_add_66132[14:11] ^ p38_add_66132[31:28], p38_add_66132[31:21] ^ p38_add_66132[10:0] ^ p38_add_66132[27:17], p38_add_66132[20:7] ^ p38_add_66132[31:18] ^ p38_add_66132[16:3]} + p38_add_65029;
  assign p39_add_67352_comb = p38_add_65844 + p39_add_67351_comb;
  assign p39_add_67333_comb = {p39_add_67306_comb[5:0] ^ p39_add_67306_comb[10:5] ^ p39_add_67306_comb[24:19], p39_add_67306_comb[31:27] ^ p39_add_67306_comb[4:0] ^ p39_add_67306_comb[18:14], p39_add_67306_comb[26:13] ^ p39_add_67306_comb[31:18] ^ p39_add_67306_comb[13:0], p39_add_67306_comb[12:6] ^ p39_add_67306_comb[17:11] ^ p39_add_67306_comb[31:25]} + p38_add_66953;
  assign p39_add_67334_comb = (p39_add_67306_comb & p38_add_67202 ^ ~(p39_add_67306_comb | ~p38_add_67102)) + {p39_add_67328_comb, p38_add_66476[1:0]};

  // Registers for pipe stage 39:
  reg [31:0] p39_add_67202;
  reg [31:0] p39_add_67306;
  reg [31:0] p39_add_66975;
  reg [31:0] p39_add_67349;
  reg [31:0] p39_add_67148;
  reg [31:0] p39_add_67252;
  reg [31:0] p39_and_67369;
  reg [31:0] p39_add_67374;
  reg [31:0] p39_add_67408;
  reg [31:0] p39_add_67391;
  reg [31:0] p39_add_66528;
  reg [31:0] p39_add_66511;
  reg [31:0] p39_add_66359;
  reg [31:0] p39_add_66624;
  reg [31:0] p39_add_66184;
  reg [31:0] p39_add_66494;
  reg [31:0] p39_add_66017;
  reg [31:0] p39_add_66325;
  reg [31:0] p39_add_67352;
  reg [31:0] p39_add_66150;
  reg [31:0] p39_add_67333;
  reg [31:0] p39_add_67334;
  reg [31:0] p39_add_66476;
  reg [31:0] p39_add_65983;
  reg [31:0] p39_add_66307;
  reg [31:0] p39_add_65810;
  always_ff @ (posedge clk) begin
    p39_add_67202 <= p38_add_67202;
    p39_add_67306 <= p39_add_67306_comb;
    p39_add_66975 <= p38_add_66975;
    p39_add_67349 <= p39_add_67349_comb;
    p39_add_67148 <= p38_add_67148;
    p39_add_67252 <= p38_add_67252;
    p39_and_67369 <= p39_and_67369_comb;
    p39_add_67374 <= p39_add_67374_comb;
    p39_add_67408 <= p39_add_67408_comb;
    p39_add_67391 <= p39_add_67391_comb;
    p39_add_66528 <= p38_add_66528;
    p39_add_66511 <= p38_add_66511;
    p39_add_66359 <= p38_add_66359;
    p39_add_66624 <= p38_add_66624;
    p39_add_66184 <= p38_add_66184;
    p39_add_66494 <= p38_add_66494;
    p39_add_66017 <= p38_add_66017;
    p39_add_66325 <= p38_add_66325;
    p39_add_67352 <= p39_add_67352_comb;
    p39_add_66150 <= p38_add_66150;
    p39_add_67333 <= p39_add_67333_comb;
    p39_add_67334 <= p39_add_67334_comb;
    p39_add_66476 <= p38_add_66476;
    p39_add_65983 <= p38_add_65983;
    p39_add_66307 <= p38_add_66307;
    p39_add_65810 <= p38_add_65810;
  end

  // ===== Pipe stage 40:
  wire [31:0] p40_add_67461_comb;
  wire [31:0] p40_add_67462_comb;
  wire [31:0] p40_and_67501_comb;
  wire [31:0] p40_add_67505_comb;
  wire [31:0] p40_add_67523_comb;
  wire [31:0] p40_add_67484_comb;
  wire [31:0] p40_add_67506_comb;
  wire [31:0] p40_add_67524_comb;
  assign p40_add_67461_comb = p39_add_67333 + p39_add_67334;
  assign p40_add_67462_comb = p39_add_66975 + p40_add_67461_comb;
  assign p40_and_67501_comb = p39_add_67374 & p39_add_67252;
  assign p40_add_67505_comb = {p39_add_67374[1:0] ^ p39_add_67374[12:11] ^ p39_add_67374[21:20], p39_add_67374[31:21] ^ p39_add_67374[10:0] ^ p39_add_67374[19:9], p39_add_67374[20:12] ^ p39_add_67374[31:23] ^ p39_add_67374[8:0], p39_add_67374[11:2] ^ p39_add_67374[22:13] ^ p39_add_67374[31:22]} + (p40_and_67501_comb ^ p39_add_67374 & p39_add_67148 ^ p39_and_67369);
  assign p40_add_67523_comb = p39_add_67352 + {p39_add_66624[16:7] ^ p39_add_66624[18:9], p39_add_66624[6:0] ^ p39_add_66624[8:2] ^ p39_add_66624[31:25], p39_add_66624[31:30] ^ p39_add_66624[1:0] ^ p39_add_66624[24:23], p39_add_66624[29:17] ^ p39_add_66624[31:19] ^ p39_add_66624[22:10]};
  assign p40_add_67484_comb = {p40_add_67462_comb[5:0] ^ p40_add_67462_comb[10:5] ^ p40_add_67462_comb[24:19], p40_add_67462_comb[31:27] ^ p40_add_67462_comb[4:0] ^ p40_add_67462_comb[18:14], p40_add_67462_comb[26:13] ^ p40_add_67462_comb[31:18] ^ p40_add_67462_comb[13:0], p40_add_67462_comb[12:6] ^ p40_add_67462_comb[17:11] ^ p40_add_67462_comb[31:25]} + (p40_add_67462_comb & p39_add_67306 ^ ~(p40_add_67462_comb | ~p39_add_67202));
  assign p40_add_67506_comb = p40_add_67461_comb + p40_add_67505_comb;
  assign p40_add_67524_comb = p39_add_66511 + p40_add_67523_comb;

  // Registers for pipe stage 40:
  reg [31:0] p40_add_67202;
  reg [31:0] p40_add_67306;
  reg [31:0] p40_add_67462;
  reg [31:0] p40_add_67484;
  reg [31:0] p40_add_67349;
  reg [31:0] p40_add_67148;
  reg [31:0] p40_add_67252;
  reg [31:0] p40_add_67374;
  reg [31:0] p40_and_67501;
  reg [31:0] p40_add_67506;
  reg [31:0] p40_add_67408;
  reg [31:0] p40_add_67391;
  reg [31:0] p40_add_66528;
  reg [31:0] p40_add_67524;
  reg [31:0] p40_add_66359;
  reg [31:0] p40_add_66624;
  reg [31:0] p40_add_66184;
  reg [31:0] p40_add_66494;
  reg [31:0] p40_add_66017;
  reg [31:0] p40_add_66325;
  reg [31:0] p40_add_67352;
  reg [31:0] p40_add_66150;
  reg [31:0] p40_add_66476;
  reg [31:0] p40_add_65983;
  reg [31:0] p40_add_66307;
  reg [31:0] p40_add_65810;
  always_ff @ (posedge clk) begin
    p40_add_67202 <= p39_add_67202;
    p40_add_67306 <= p39_add_67306;
    p40_add_67462 <= p40_add_67462_comb;
    p40_add_67484 <= p40_add_67484_comb;
    p40_add_67349 <= p39_add_67349;
    p40_add_67148 <= p39_add_67148;
    p40_add_67252 <= p39_add_67252;
    p40_add_67374 <= p39_add_67374;
    p40_and_67501 <= p40_and_67501_comb;
    p40_add_67506 <= p40_add_67506_comb;
    p40_add_67408 <= p39_add_67408;
    p40_add_67391 <= p39_add_67391;
    p40_add_66528 <= p39_add_66528;
    p40_add_67524 <= p40_add_67524_comb;
    p40_add_66359 <= p39_add_66359;
    p40_add_66624 <= p39_add_66624;
    p40_add_66184 <= p39_add_66184;
    p40_add_66494 <= p39_add_66494;
    p40_add_66017 <= p39_add_66017;
    p40_add_66325 <= p39_add_66325;
    p40_add_67352 <= p39_add_67352;
    p40_add_66150 <= p39_add_66150;
    p40_add_66476 <= p39_add_66476;
    p40_add_65983 <= p39_add_65983;
    p40_add_66307 <= p39_add_66307;
    p40_add_65810 <= p39_add_65810;
  end

  // ===== Pipe stage 41:
  wire [31:0] p41_and_67600_comb;
  wire [31:0] p41_add_67578_comb;
  wire [31:0] p41_add_67579_comb;
  wire [31:0] p41_add_67604_comb;
  wire [31:0] p41_add_67580_comb;
  wire [29:0] p41_add_67583_comb;
  wire [31:0] p41_add_67605_comb;
  assign p41_and_67600_comb = p40_add_67506 & p40_add_67374;
  assign p41_add_67578_comb = p40_add_67484 + 32'h5338_0d13;
  assign p41_add_67579_comb = p41_add_67578_comb + p40_add_67349;
  assign p41_add_67604_comb = {p40_add_67506[1:0] ^ p40_add_67506[12:11] ^ p40_add_67506[21:20], p40_add_67506[31:21] ^ p40_add_67506[10:0] ^ p40_add_67506[19:9], p40_add_67506[20:12] ^ p40_add_67506[31:23] ^ p40_add_67506[8:0], p40_add_67506[11:2] ^ p40_add_67506[22:13] ^ p40_add_67506[31:22]} + (p41_and_67600_comb ^ p40_add_67506 & p40_add_67252 ^ p40_and_67501);
  assign p41_add_67580_comb = p40_add_67148 + p41_add_67579_comb;
  assign p41_add_67583_comb = p40_add_67352[31:2] + 30'h1942_9cd5;
  assign p41_add_67605_comb = p41_add_67579_comb + p41_add_67604_comb;

  // Registers for pipe stage 41:
  reg [31:0] p41_add_67202;
  reg [31:0] p41_add_67306;
  reg [31:0] p41_add_67462;
  reg [31:0] p41_add_67580;
  reg [29:0] p41_add_67583;
  reg [31:0] p41_add_67252;
  reg [31:0] p41_add_67374;
  reg [31:0] p41_add_67506;
  reg [31:0] p41_and_67600;
  reg [31:0] p41_add_67605;
  reg [31:0] p41_add_67408;
  reg [31:0] p41_add_67391;
  reg [31:0] p41_add_66528;
  reg [31:0] p41_add_67524;
  reg [31:0] p41_add_66359;
  reg [31:0] p41_add_66624;
  reg [31:0] p41_add_66184;
  reg [31:0] p41_add_66494;
  reg [31:0] p41_add_66017;
  reg [31:0] p41_add_66325;
  reg [31:0] p41_add_67352;
  reg [31:0] p41_add_66150;
  reg [31:0] p41_add_66476;
  reg [31:0] p41_add_65983;
  reg [31:0] p41_add_66307;
  reg [31:0] p41_add_65810;
  always_ff @ (posedge clk) begin
    p41_add_67202 <= p40_add_67202;
    p41_add_67306 <= p40_add_67306;
    p41_add_67462 <= p40_add_67462;
    p41_add_67580 <= p41_add_67580_comb;
    p41_add_67583 <= p41_add_67583_comb;
    p41_add_67252 <= p40_add_67252;
    p41_add_67374 <= p40_add_67374;
    p41_add_67506 <= p40_add_67506;
    p41_and_67600 <= p41_and_67600_comb;
    p41_add_67605 <= p41_add_67605_comb;
    p41_add_67408 <= p40_add_67408;
    p41_add_67391 <= p40_add_67391;
    p41_add_66528 <= p40_add_66528;
    p41_add_67524 <= p40_add_67524;
    p41_add_66359 <= p40_add_66359;
    p41_add_66624 <= p40_add_66624;
    p41_add_66184 <= p40_add_66184;
    p41_add_66494 <= p40_add_66494;
    p41_add_66017 <= p40_add_66017;
    p41_add_66325 <= p40_add_66325;
    p41_add_67352 <= p40_add_67352;
    p41_add_66150 <= p40_add_66150;
    p41_add_66476 <= p40_add_66476;
    p41_add_65983 <= p40_add_65983;
    p41_add_66307 <= p40_add_66307;
    p41_add_65810 <= p40_add_65810;
  end

  // ===== Pipe stage 42:
  wire [31:0] p42_and_67719_comb;
  wire [31:0] p42_add_67681_comb;
  wire [31:0] p42_add_67682_comb;
  wire [31:0] p42_add_67683_comb;
  wire [31:0] p42_add_67723_comb;
  wire [31:0] p42_add_67701_comb;
  wire [31:0] p42_add_67684_comb;
  wire [31:0] p42_add_67699_comb;
  wire [31:0] p42_add_67724_comb;
  wire [31:0] p42_add_67758_comb;
  wire [31:0] p42_add_67741_comb;
  wire [31:0] p42_add_67702_comb;
  assign p42_and_67719_comb = p41_add_67605 & p41_add_67506;
  assign p42_add_67681_comb = {p41_add_67580[5:0] ^ p41_add_67580[10:5] ^ p41_add_67580[24:19], p41_add_67580[31:27] ^ p41_add_67580[4:0] ^ p41_add_67580[18:14], p41_add_67580[26:13] ^ p41_add_67580[31:18] ^ p41_add_67580[13:0], p41_add_67580[12:6] ^ p41_add_67580[17:11] ^ p41_add_67580[31:25]} + p41_add_67202;
  assign p42_add_67682_comb = (p41_add_67580 & p41_add_67462 ^ ~(p41_add_67580 | ~p41_add_67306)) + {p41_add_67583, p41_add_67352[1:0]};
  assign p42_add_67683_comb = p42_add_67681_comb + p42_add_67682_comb;
  assign p42_add_67723_comb = {p41_add_67605[1:0] ^ p41_add_67605[12:11] ^ p41_add_67605[21:20], p41_add_67605[31:21] ^ p41_add_67605[10:0] ^ p41_add_67605[19:9], p41_add_67605[20:12] ^ p41_add_67605[31:23] ^ p41_add_67605[8:0], p41_add_67605[11:2] ^ p41_add_67605[22:13] ^ p41_add_67605[31:22]} + (p42_and_67719_comb ^ p41_add_67605 & p41_add_67374 ^ p41_and_67600);
  assign p42_add_67701_comb = p41_add_65810 + {p41_add_67352[16:7] ^ p41_add_67352[18:9], p41_add_67352[6:0] ^ p41_add_67352[8:2] ^ p41_add_67352[31:25], p41_add_67352[31:30] ^ p41_add_67352[1:0] ^ p41_add_67352[24:23], p41_add_67352[29:17] ^ p41_add_67352[31:19] ^ p41_add_67352[22:10]};
  assign p42_add_67684_comb = p41_add_67252 + p42_add_67683_comb;
  assign p42_add_67699_comb = p41_add_67306 + p41_add_66325;
  assign p42_add_67724_comb = p42_add_67683_comb + p42_add_67723_comb;
  assign p42_add_67758_comb = {p41_add_65983[6:4] ^ p41_add_65983[17:15], p41_add_65983[3:0] ^ p41_add_65983[14:11] ^ p41_add_65983[31:28], p41_add_65983[31:21] ^ p41_add_65983[10:0] ^ p41_add_65983[27:17], p41_add_65983[20:7] ^ p41_add_65983[31:18] ^ p41_add_65983[16:3]} + p41_add_66307;
  assign p42_add_67741_comb = {p41_add_66307[6:4] ^ p41_add_66307[17:15], p41_add_66307[3:0] ^ p41_add_66307[14:11] ^ p41_add_66307[31:28], p41_add_66307[31:21] ^ p41_add_66307[10:0] ^ p41_add_66307[27:17], p41_add_66307[20:7] ^ p41_add_66307[31:18] ^ p41_add_66307[16:3]} + p41_add_65810;
  assign p42_add_67702_comb = p41_add_66017 + p42_add_67701_comb;

  // Registers for pipe stage 42:
  reg [31:0] p42_add_67462;
  reg [31:0] p42_add_67580;
  reg [31:0] p42_add_67684;
  reg [31:0] p42_add_67699;
  reg [31:0] p42_add_67374;
  reg [31:0] p42_add_67506;
  reg [31:0] p42_add_67605;
  reg [31:0] p42_and_67719;
  reg [31:0] p42_add_67724;
  reg [31:0] p42_add_67758;
  reg [31:0] p42_add_67741;
  reg [31:0] p42_add_67408;
  reg [31:0] p42_add_67391;
  reg [31:0] p42_add_66528;
  reg [31:0] p42_add_67524;
  reg [31:0] p42_add_66359;
  reg [31:0] p42_add_66624;
  reg [31:0] p42_add_66184;
  reg [31:0] p42_add_66494;
  reg [31:0] p42_add_67702;
  reg [31:0] p42_add_66325;
  reg [31:0] p42_add_67352;
  reg [31:0] p42_add_66150;
  reg [31:0] p42_add_66476;
  reg [31:0] p42_add_65983;
  always_ff @ (posedge clk) begin
    p42_add_67462 <= p41_add_67462;
    p42_add_67580 <= p41_add_67580;
    p42_add_67684 <= p42_add_67684_comb;
    p42_add_67699 <= p42_add_67699_comb;
    p42_add_67374 <= p41_add_67374;
    p42_add_67506 <= p41_add_67506;
    p42_add_67605 <= p41_add_67605;
    p42_and_67719 <= p42_and_67719_comb;
    p42_add_67724 <= p42_add_67724_comb;
    p42_add_67758 <= p42_add_67758_comb;
    p42_add_67741 <= p42_add_67741_comb;
    p42_add_67408 <= p41_add_67408;
    p42_add_67391 <= p41_add_67391;
    p42_add_66528 <= p41_add_66528;
    p42_add_67524 <= p41_add_67524;
    p42_add_66359 <= p41_add_66359;
    p42_add_66624 <= p41_add_66624;
    p42_add_66184 <= p41_add_66184;
    p42_add_66494 <= p41_add_66494;
    p42_add_67702 <= p42_add_67702_comb;
    p42_add_66325 <= p41_add_66325;
    p42_add_67352 <= p41_add_67352;
    p42_add_66150 <= p41_add_66150;
    p42_add_66476 <= p41_add_66476;
    p42_add_65983 <= p41_add_65983;
  end

  // ===== Pipe stage 43:
  wire [31:0] p43_add_67830_comb;
  wire [31:0] p43_add_67832_comb;
  wire [31:0] p43_add_67868_comb;
  wire [31:0] p43_add_67850_comb;
  wire [31:0] p43_add_67833_comb;
  wire [31:0] p43_add_67903_comb;
  wire [31:0] p43_add_67886_comb;
  wire [31:0] p43_add_67869_comb;
  wire [31:0] p43_add_67851_comb;
  assign p43_add_67830_comb = {p42_add_67684[5:0] ^ p42_add_67684[10:5] ^ p42_add_67684[24:19], p42_add_67684[31:27] ^ p42_add_67684[4:0] ^ p42_add_67684[18:14], p42_add_67684[26:13] ^ p42_add_67684[31:18] ^ p42_add_67684[13:0], p42_add_67684[12:6] ^ p42_add_67684[17:11] ^ p42_add_67684[31:25]} + (p42_add_67684 & p42_add_67580 ^ ~(p42_add_67684 | ~p42_add_67462));
  assign p43_add_67832_comb = p43_add_67830_comb + 32'h766a_0abb;
  assign p43_add_67868_comb = p42_add_67702 + {p42_add_67524[16:7] ^ p42_add_67524[18:9], p42_add_67524[6:0] ^ p42_add_67524[8:2] ^ p42_add_67524[31:25], p42_add_67524[31:30] ^ p42_add_67524[1:0] ^ p42_add_67524[24:23], p42_add_67524[29:17] ^ p42_add_67524[31:19] ^ p42_add_67524[22:10]};
  assign p43_add_67850_comb = p42_add_65983 + {p42_add_67702[16:7] ^ p42_add_67702[18:9], p42_add_67702[6:0] ^ p42_add_67702[8:2] ^ p42_add_67702[31:25], p42_add_67702[31:30] ^ p42_add_67702[1:0] ^ p42_add_67702[24:23], p42_add_67702[29:17] ^ p42_add_67702[31:19] ^ p42_add_67702[22:10]};
  assign p43_add_67833_comb = p43_add_67832_comb + p42_add_67699;
  assign p43_add_67903_comb = {p42_add_66150[6:4] ^ p42_add_66150[17:15], p42_add_66150[3:0] ^ p42_add_66150[14:11] ^ p42_add_66150[31:28], p42_add_66150[31:21] ^ p42_add_66150[10:0] ^ p42_add_66150[27:17], p42_add_66150[20:7] ^ p42_add_66150[31:18] ^ p42_add_66150[16:3]} + p42_add_66476;
  assign p43_add_67886_comb = {p42_add_66476[6:4] ^ p42_add_66476[17:15], p42_add_66476[3:0] ^ p42_add_66476[14:11] ^ p42_add_66476[31:28], p42_add_66476[31:21] ^ p42_add_66476[10:0] ^ p42_add_66476[27:17], p42_add_66476[20:7] ^ p42_add_66476[31:18] ^ p42_add_66476[16:3]} + p42_add_65983;
  assign p43_add_67869_comb = p42_add_67391 + p43_add_67868_comb;
  assign p43_add_67851_comb = p42_add_66184 + p43_add_67850_comb;

  // Registers for pipe stage 43:
  reg [31:0] p43_add_67462;
  reg [31:0] p43_add_67580;
  reg [31:0] p43_add_67684;
  reg [31:0] p43_add_67374;
  reg [31:0] p43_add_67833;
  reg [31:0] p43_add_67506;
  reg [31:0] p43_add_67605;
  reg [31:0] p43_and_67719;
  reg [31:0] p43_add_67724;
  reg [31:0] p43_add_67903;
  reg [31:0] p43_add_67886;
  reg [31:0] p43_add_67758;
  reg [31:0] p43_add_67741;
  reg [31:0] p43_add_67408;
  reg [31:0] p43_add_67869;
  reg [31:0] p43_add_66528;
  reg [31:0] p43_add_67524;
  reg [31:0] p43_add_66359;
  reg [31:0] p43_add_66624;
  reg [31:0] p43_add_67851;
  reg [31:0] p43_add_66494;
  reg [31:0] p43_add_67702;
  reg [31:0] p43_add_66325;
  reg [31:0] p43_add_67352;
  reg [31:0] p43_add_66150;
  always_ff @ (posedge clk) begin
    p43_add_67462 <= p42_add_67462;
    p43_add_67580 <= p42_add_67580;
    p43_add_67684 <= p42_add_67684;
    p43_add_67374 <= p42_add_67374;
    p43_add_67833 <= p43_add_67833_comb;
    p43_add_67506 <= p42_add_67506;
    p43_add_67605 <= p42_add_67605;
    p43_and_67719 <= p42_and_67719;
    p43_add_67724 <= p42_add_67724;
    p43_add_67903 <= p43_add_67903_comb;
    p43_add_67886 <= p43_add_67886_comb;
    p43_add_67758 <= p42_add_67758;
    p43_add_67741 <= p42_add_67741;
    p43_add_67408 <= p42_add_67408;
    p43_add_67869 <= p43_add_67869_comb;
    p43_add_66528 <= p42_add_66528;
    p43_add_67524 <= p42_add_67524;
    p43_add_66359 <= p42_add_66359;
    p43_add_66624 <= p42_add_66624;
    p43_add_67851 <= p43_add_67851_comb;
    p43_add_66494 <= p42_add_66494;
    p43_add_67702 <= p42_add_67702;
    p43_add_66325 <= p42_add_66325;
    p43_add_67352 <= p42_add_67352;
    p43_add_66150 <= p42_add_66150;
  end

  // ===== Pipe stage 44:
  wire [31:0] p44_add_67954_comb;
  wire [31:0] p44_and_68001_comb;
  wire [30:0] p44_add_67976_comb;
  wire [31:0] p44_add_68020_comb;
  wire [31:0] p44_add_68023_comb;
  wire [31:0] p44_add_67981_comb;
  wire [31:0] p44_add_67982_comb;
  wire [31:0] p44_add_67984_comb;
  wire [31:0] p44_add_68022_comb;
  wire [31:0] p44_add_68058_comb;
  wire [31:0] p44_add_68041_comb;
  wire [31:0] p44_add_68024_comb;
  wire [31:0] p44_add_67983_comb;
  assign p44_add_67954_comb = p43_add_67374 + p43_add_67833;
  assign p44_and_68001_comb = p43_add_67724 & p43_add_67605;
  assign p44_add_67976_comb = p43_add_67702[31:1] + 31'h40e1_6497;
  assign p44_add_68020_comb = {p43_add_67724[1:0] ^ p43_add_67724[12:11] ^ p43_add_67724[21:20], p43_add_67724[31:21] ^ p43_add_67724[10:0] ^ p43_add_67724[19:9], p43_add_67724[20:12] ^ p43_add_67724[31:23] ^ p43_add_67724[8:0], p43_add_67724[11:2] ^ p43_add_67724[22:13] ^ p43_add_67724[31:22]} + (p44_and_68001_comb ^ p43_add_67724 & p43_add_67506 ^ p43_and_67719);
  assign p44_add_68023_comb = p43_add_66150 + {p43_add_67851[16:7] ^ p43_add_67851[18:9], p43_add_67851[6:0] ^ p43_add_67851[8:2] ^ p43_add_67851[31:25], p43_add_67851[31:30] ^ p43_add_67851[1:0] ^ p43_add_67851[24:23], p43_add_67851[29:17] ^ p43_add_67851[31:19] ^ p43_add_67851[22:10]};
  assign p44_add_67981_comb = {p44_add_67954_comb[5:0] ^ p44_add_67954_comb[10:5] ^ p44_add_67954_comb[24:19], p44_add_67954_comb[31:27] ^ p44_add_67954_comb[4:0] ^ p44_add_67954_comb[18:14], p44_add_67954_comb[26:13] ^ p44_add_67954_comb[31:18] ^ p44_add_67954_comb[13:0], p44_add_67954_comb[12:6] ^ p44_add_67954_comb[17:11] ^ p44_add_67954_comb[31:25]} + p43_add_67462;
  assign p44_add_67982_comb = (p44_add_67954_comb & p43_add_67684 ^ ~(p44_add_67954_comb | ~p43_add_67580)) + {p44_add_67976_comb, p43_add_67702[0]};
  assign p44_add_67984_comb = p43_add_67580 + p43_add_66494;
  assign p44_add_68022_comb = p43_add_67833 + p44_add_68020_comb;
  assign p44_add_68058_comb = {p43_add_66325[6:4] ^ p43_add_66325[17:15], p43_add_66325[3:0] ^ p43_add_66325[14:11] ^ p43_add_66325[31:28], p43_add_66325[31:21] ^ p43_add_66325[10:0] ^ p43_add_66325[27:17], p43_add_66325[20:7] ^ p43_add_66325[31:18] ^ p43_add_66325[16:3]} + p43_add_67352;
  assign p44_add_68041_comb = {p43_add_67352[6:4] ^ p43_add_67352[17:15], p43_add_67352[3:0] ^ p43_add_67352[14:11] ^ p43_add_67352[31:28], p43_add_67352[31:21] ^ p43_add_67352[10:0] ^ p43_add_67352[27:17], p43_add_67352[20:7] ^ p43_add_67352[31:18] ^ p43_add_67352[16:3]} + p43_add_66150;
  assign p44_add_68024_comb = p43_add_66359 + p44_add_68023_comb;
  assign p44_add_67983_comb = p44_add_67981_comb + p44_add_67982_comb;

  // Registers for pipe stage 44:
  reg [31:0] p44_add_67684;
  reg [31:0] p44_add_67954;
  reg [31:0] p44_add_67506;
  reg [31:0] p44_add_67984;
  reg [31:0] p44_add_67605;
  reg [31:0] p44_add_67724;
  reg [31:0] p44_and_68001;
  reg [31:0] p44_add_68022;
  reg [31:0] p44_add_68058;
  reg [31:0] p44_add_68041;
  reg [31:0] p44_add_67903;
  reg [31:0] p44_add_67886;
  reg [31:0] p44_add_67758;
  reg [31:0] p44_add_67741;
  reg [31:0] p44_add_67408;
  reg [31:0] p44_add_67869;
  reg [31:0] p44_add_66528;
  reg [31:0] p44_add_67524;
  reg [31:0] p44_add_68024;
  reg [31:0] p44_add_66624;
  reg [31:0] p44_add_67851;
  reg [31:0] p44_add_66494;
  reg [31:0] p44_add_67983;
  reg [31:0] p44_add_67702;
  reg [31:0] p44_add_66325;
  always_ff @ (posedge clk) begin
    p44_add_67684 <= p43_add_67684;
    p44_add_67954 <= p44_add_67954_comb;
    p44_add_67506 <= p43_add_67506;
    p44_add_67984 <= p44_add_67984_comb;
    p44_add_67605 <= p43_add_67605;
    p44_add_67724 <= p43_add_67724;
    p44_and_68001 <= p44_and_68001_comb;
    p44_add_68022 <= p44_add_68022_comb;
    p44_add_68058 <= p44_add_68058_comb;
    p44_add_68041 <= p44_add_68041_comb;
    p44_add_67903 <= p43_add_67903;
    p44_add_67886 <= p43_add_67886;
    p44_add_67758 <= p43_add_67758;
    p44_add_67741 <= p43_add_67741;
    p44_add_67408 <= p43_add_67408;
    p44_add_67869 <= p43_add_67869;
    p44_add_66528 <= p43_add_66528;
    p44_add_67524 <= p43_add_67524;
    p44_add_68024 <= p44_add_68024_comb;
    p44_add_66624 <= p43_add_66624;
    p44_add_67851 <= p43_add_67851;
    p44_add_66494 <= p43_add_66494;
    p44_add_67983 <= p44_add_67983_comb;
    p44_add_67702 <= p43_add_67702;
    p44_add_66325 <= p43_add_66325;
  end

  // ===== Pipe stage 45:
  wire [31:0] p45_add_68109_comb;
  wire [31:0] p45_and_68151_comb;
  wire [31:0] p45_add_68155_comb;
  wire [31:0] p45_add_68131_comb;
  wire [31:0] p45_add_68173_comb;
  wire [31:0] p45_add_68134_comb;
  wire [31:0] p45_add_68156_comb;
  wire [31:0] p45_add_68133_comb;
  wire [31:0] p45_add_68208_comb;
  wire [31:0] p45_add_68191_comb;
  wire [31:0] p45_add_68174_comb;
  assign p45_add_68109_comb = p44_add_67506 + p44_add_67983;
  assign p45_and_68151_comb = p44_add_68022 & p44_add_67724;
  assign p45_add_68155_comb = {p44_add_68022[1:0] ^ p44_add_68022[12:11] ^ p44_add_68022[21:20], p44_add_68022[31:21] ^ p44_add_68022[10:0] ^ p44_add_68022[19:9], p44_add_68022[20:12] ^ p44_add_68022[31:23] ^ p44_add_68022[8:0], p44_add_68022[11:2] ^ p44_add_68022[22:13] ^ p44_add_68022[31:22]} + (p45_and_68151_comb ^ p44_add_68022 & p44_add_67605 ^ p44_and_68001);
  assign p45_add_68131_comb = {p45_add_68109_comb[5:0] ^ p45_add_68109_comb[10:5] ^ p45_add_68109_comb[24:19], p45_add_68109_comb[31:27] ^ p45_add_68109_comb[4:0] ^ p45_add_68109_comb[18:14], p45_add_68109_comb[26:13] ^ p45_add_68109_comb[31:18] ^ p45_add_68109_comb[13:0], p45_add_68109_comb[12:6] ^ p45_add_68109_comb[17:11] ^ p45_add_68109_comb[31:25]} + (p45_add_68109_comb & p44_add_67954 ^ ~(p45_add_68109_comb | ~p44_add_67684));
  assign p45_add_68173_comb = p44_add_66325 + {p44_add_68024[16:7] ^ p44_add_68024[18:9], p44_add_68024[6:0] ^ p44_add_68024[8:2] ^ p44_add_68024[31:25], p44_add_68024[31:30] ^ p44_add_68024[1:0] ^ p44_add_68024[24:23], p44_add_68024[29:17] ^ p44_add_68024[31:19] ^ p44_add_68024[22:10]};
  assign p45_add_68134_comb = p44_add_67684 + p44_add_67851;
  assign p45_add_68156_comb = p44_add_67983 + p45_add_68155_comb;
  assign p45_add_68133_comb = p45_add_68131_comb + 32'h9272_2c85;
  assign p45_add_68208_comb = {p44_add_66494[6:4] ^ p44_add_66494[17:15], p44_add_66494[3:0] ^ p44_add_66494[14:11] ^ p44_add_66494[31:28], p44_add_66494[31:21] ^ p44_add_66494[10:0] ^ p44_add_66494[27:17], p44_add_66494[20:7] ^ p44_add_66494[31:18] ^ p44_add_66494[16:3]} + p44_add_67702;
  assign p45_add_68191_comb = {p44_add_67702[6:4] ^ p44_add_67702[17:15], p44_add_67702[3:0] ^ p44_add_67702[14:11] ^ p44_add_67702[31:28], p44_add_67702[31:21] ^ p44_add_67702[10:0] ^ p44_add_67702[27:17], p44_add_67702[20:7] ^ p44_add_67702[31:18] ^ p44_add_67702[16:3]} + p44_add_66325;
  assign p45_add_68174_comb = p44_add_66528 + p45_add_68173_comb;

  // Registers for pipe stage 45:
  reg [31:0] p45_add_67954;
  reg [31:0] p45_add_68109;
  reg [31:0] p45_add_67984;
  reg [31:0] p45_add_67605;
  reg [31:0] p45_add_68134;
  reg [31:0] p45_add_67724;
  reg [31:0] p45_add_68022;
  reg [31:0] p45_and_68151;
  reg [31:0] p45_add_68156;
  reg [31:0] p45_add_68133;
  reg [31:0] p45_add_68208;
  reg [31:0] p45_add_68191;
  reg [31:0] p45_add_68058;
  reg [31:0] p45_add_68041;
  reg [31:0] p45_add_67903;
  reg [31:0] p45_add_67886;
  reg [31:0] p45_add_67758;
  reg [31:0] p45_add_67741;
  reg [31:0] p45_add_67408;
  reg [31:0] p45_add_67869;
  reg [31:0] p45_add_68174;
  reg [31:0] p45_add_67524;
  reg [31:0] p45_add_68024;
  reg [31:0] p45_add_66624;
  reg [31:0] p45_add_67851;
  reg [31:0] p45_add_66494;
  always_ff @ (posedge clk) begin
    p45_add_67954 <= p44_add_67954;
    p45_add_68109 <= p45_add_68109_comb;
    p45_add_67984 <= p44_add_67984;
    p45_add_67605 <= p44_add_67605;
    p45_add_68134 <= p45_add_68134_comb;
    p45_add_67724 <= p44_add_67724;
    p45_add_68022 <= p44_add_68022;
    p45_and_68151 <= p45_and_68151_comb;
    p45_add_68156 <= p45_add_68156_comb;
    p45_add_68133 <= p45_add_68133_comb;
    p45_add_68208 <= p45_add_68208_comb;
    p45_add_68191 <= p45_add_68191_comb;
    p45_add_68058 <= p44_add_68058;
    p45_add_68041 <= p44_add_68041;
    p45_add_67903 <= p44_add_67903;
    p45_add_67886 <= p44_add_67886;
    p45_add_67758 <= p44_add_67758;
    p45_add_67741 <= p44_add_67741;
    p45_add_67408 <= p44_add_67408;
    p45_add_67869 <= p44_add_67869;
    p45_add_68174 <= p45_add_68174_comb;
    p45_add_67524 <= p44_add_67524;
    p45_add_68024 <= p44_add_68024;
    p45_add_66624 <= p44_add_66624;
    p45_add_67851 <= p44_add_67851;
    p45_add_66494 <= p44_add_66494;
  end

  // ===== Pipe stage 46:
  wire [31:0] p46_add_68261_comb;
  wire [31:0] p46_add_68262_comb;
  wire [31:0] p46_and_68302_comb;
  wire [31:0] p46_add_68306_comb;
  wire [31:0] p46_add_68324_comb;
  wire [31:0] p46_add_68284_comb;
  wire [31:0] p46_add_68285_comb;
  wire [31:0] p46_add_68307_comb;
  wire [31:0] p46_add_68342_comb;
  wire [31:0] p46_add_68325_comb;
  assign p46_add_68261_comb = p45_add_68133 + p45_add_67984;
  assign p46_add_68262_comb = p45_add_67605 + p46_add_68261_comb;
  assign p46_and_68302_comb = p45_add_68156 & p45_add_68022;
  assign p46_add_68306_comb = {p45_add_68156[1:0] ^ p45_add_68156[12:11] ^ p45_add_68156[21:20], p45_add_68156[31:21] ^ p45_add_68156[10:0] ^ p45_add_68156[19:9], p45_add_68156[20:12] ^ p45_add_68156[31:23] ^ p45_add_68156[8:0], p45_add_68156[11:2] ^ p45_add_68156[22:13] ^ p45_add_68156[31:22]} + (p46_and_68302_comb ^ p45_add_68156 & p45_add_67724 ^ p45_and_68151);
  assign p46_add_68324_comb = p45_add_66494 + {p45_add_68174[16:7] ^ p45_add_68174[18:9], p45_add_68174[6:0] ^ p45_add_68174[8:2] ^ p45_add_68174[31:25], p45_add_68174[31:30] ^ p45_add_68174[1:0] ^ p45_add_68174[24:23], p45_add_68174[29:17] ^ p45_add_68174[31:19] ^ p45_add_68174[22:10]};
  assign p46_add_68284_comb = {p46_add_68262_comb[5:0] ^ p46_add_68262_comb[10:5] ^ p46_add_68262_comb[24:19], p46_add_68262_comb[31:27] ^ p46_add_68262_comb[4:0] ^ p46_add_68262_comb[18:14], p46_add_68262_comb[26:13] ^ p46_add_68262_comb[31:18] ^ p46_add_68262_comb[13:0], p46_add_68262_comb[12:6] ^ p46_add_68262_comb[17:11] ^ p46_add_68262_comb[31:25]} + (p46_add_68262_comb & p45_add_68109 ^ ~(p46_add_68262_comb | ~p45_add_67954));
  assign p46_add_68285_comb = p45_add_67954 + p45_add_66624;
  assign p46_add_68307_comb = p46_add_68261_comb + p46_add_68306_comb;
  assign p46_add_68342_comb = {p45_add_67851[6:4] ^ p45_add_67851[17:15], p45_add_67851[3:0] ^ p45_add_67851[14:11] ^ p45_add_67851[31:28], p45_add_67851[31:21] ^ p45_add_67851[10:0] ^ p45_add_67851[27:17], p45_add_67851[20:7] ^ p45_add_67851[31:18] ^ p45_add_67851[16:3]} + p45_add_66494;
  assign p46_add_68325_comb = p45_add_67408 + p46_add_68324_comb;

  // Registers for pipe stage 46:
  reg [31:0] p46_add_68109;
  reg [31:0] p46_add_68262;
  reg [31:0] p46_add_68284;
  reg [31:0] p46_add_68134;
  reg [31:0] p46_add_67724;
  reg [31:0] p46_add_68285;
  reg [31:0] p46_add_68022;
  reg [31:0] p46_add_68156;
  reg [31:0] p46_and_68302;
  reg [31:0] p46_add_68307;
  reg [31:0] p46_add_68342;
  reg [31:0] p46_add_68208;
  reg [31:0] p46_add_68191;
  reg [31:0] p46_add_68058;
  reg [31:0] p46_add_68041;
  reg [31:0] p46_add_67903;
  reg [31:0] p46_add_67886;
  reg [31:0] p46_add_67758;
  reg [31:0] p46_add_67741;
  reg [31:0] p46_add_68325;
  reg [31:0] p46_add_67869;
  reg [31:0] p46_add_68174;
  reg [31:0] p46_add_67524;
  reg [31:0] p46_add_68024;
  reg [31:0] p46_add_66624;
  reg [31:0] p46_add_67851;
  always_ff @ (posedge clk) begin
    p46_add_68109 <= p45_add_68109;
    p46_add_68262 <= p46_add_68262_comb;
    p46_add_68284 <= p46_add_68284_comb;
    p46_add_68134 <= p45_add_68134;
    p46_add_67724 <= p45_add_67724;
    p46_add_68285 <= p46_add_68285_comb;
    p46_add_68022 <= p45_add_68022;
    p46_add_68156 <= p45_add_68156;
    p46_and_68302 <= p46_and_68302_comb;
    p46_add_68307 <= p46_add_68307_comb;
    p46_add_68342 <= p46_add_68342_comb;
    p46_add_68208 <= p45_add_68208;
    p46_add_68191 <= p45_add_68191;
    p46_add_68058 <= p45_add_68058;
    p46_add_68041 <= p45_add_68041;
    p46_add_67903 <= p45_add_67903;
    p46_add_67886 <= p45_add_67886;
    p46_add_67758 <= p45_add_67758;
    p46_add_67741 <= p45_add_67741;
    p46_add_68325 <= p46_add_68325_comb;
    p46_add_67869 <= p45_add_67869;
    p46_add_68174 <= p45_add_68174;
    p46_add_67524 <= p45_add_67524;
    p46_add_68024 <= p45_add_68024;
    p46_add_66624 <= p45_add_66624;
    p46_add_67851 <= p45_add_67851;
  end

  // ===== Pipe stage 47:
  wire [31:0] p47_and_68415_comb;
  wire [31:0] p47_add_68396_comb;
  wire [31:0] p47_add_68397_comb;
  wire [31:0] p47_add_68419_comb;
  wire [31:0] p47_add_68437_comb;
  wire [31:0] p47_add_68398_comb;
  wire [31:0] p47_add_68420_comb;
  wire [31:0] p47_add_68438_comb;
  assign p47_and_68415_comb = p46_add_68307 & p46_add_68156;
  assign p47_add_68396_comb = p46_add_68284 + 32'ha2bf_e8a1;
  assign p47_add_68397_comb = p47_add_68396_comb + p46_add_68134;
  assign p47_add_68419_comb = {p46_add_68307[1:0] ^ p46_add_68307[12:11] ^ p46_add_68307[21:20], p46_add_68307[31:21] ^ p46_add_68307[10:0] ^ p46_add_68307[19:9], p46_add_68307[20:12] ^ p46_add_68307[31:23] ^ p46_add_68307[8:0], p46_add_68307[11:2] ^ p46_add_68307[22:13] ^ p46_add_68307[31:22]} + (p47_and_68415_comb ^ p46_add_68307 & p46_add_68022 ^ p46_and_68302);
  assign p47_add_68437_comb = p46_add_66624 + {p46_add_68325[16:7] ^ p46_add_68325[18:9], p46_add_68325[6:0] ^ p46_add_68325[8:2] ^ p46_add_68325[31:25], p46_add_68325[31:30] ^ p46_add_68325[1:0] ^ p46_add_68325[24:23], p46_add_68325[29:17] ^ p46_add_68325[31:19] ^ p46_add_68325[22:10]};
  assign p47_add_68398_comb = p46_add_67724 + p47_add_68397_comb;
  assign p47_add_68420_comb = p47_add_68397_comb + p47_add_68419_comb;
  assign p47_add_68438_comb = p46_add_67758 + p47_add_68437_comb;

  // Registers for pipe stage 47:
  reg [31:0] p47_add_68109;
  reg [31:0] p47_add_68262;
  reg [31:0] p47_add_68398;
  reg [31:0] p47_add_68285;
  reg [31:0] p47_add_68022;
  reg [31:0] p47_add_68156;
  reg [31:0] p47_add_68307;
  reg [31:0] p47_and_68415;
  reg [31:0] p47_add_68420;
  reg [31:0] p47_add_68342;
  reg [31:0] p47_add_68208;
  reg [31:0] p47_add_68191;
  reg [31:0] p47_add_68058;
  reg [31:0] p47_add_68041;
  reg [31:0] p47_add_67903;
  reg [31:0] p47_add_67886;
  reg [31:0] p47_add_68438;
  reg [31:0] p47_add_67741;
  reg [31:0] p47_add_68325;
  reg [31:0] p47_add_67869;
  reg [31:0] p47_add_68174;
  reg [31:0] p47_add_67524;
  reg [31:0] p47_add_68024;
  reg [31:0] p47_add_66624;
  reg [31:0] p47_add_67851;
  always_ff @ (posedge clk) begin
    p47_add_68109 <= p46_add_68109;
    p47_add_68262 <= p46_add_68262;
    p47_add_68398 <= p47_add_68398_comb;
    p47_add_68285 <= p46_add_68285;
    p47_add_68022 <= p46_add_68022;
    p47_add_68156 <= p46_add_68156;
    p47_add_68307 <= p46_add_68307;
    p47_and_68415 <= p47_and_68415_comb;
    p47_add_68420 <= p47_add_68420_comb;
    p47_add_68342 <= p46_add_68342;
    p47_add_68208 <= p46_add_68208;
    p47_add_68191 <= p46_add_68191;
    p47_add_68058 <= p46_add_68058;
    p47_add_68041 <= p46_add_68041;
    p47_add_67903 <= p46_add_67903;
    p47_add_67886 <= p46_add_67886;
    p47_add_68438 <= p47_add_68438_comb;
    p47_add_67741 <= p46_add_67741;
    p47_add_68325 <= p46_add_68325;
    p47_add_67869 <= p46_add_67869;
    p47_add_68174 <= p46_add_68174;
    p47_add_67524 <= p46_add_67524;
    p47_add_68024 <= p46_add_68024;
    p47_add_66624 <= p46_add_66624;
    p47_add_67851 <= p46_add_67851;
  end

  // ===== Pipe stage 48:
  wire [31:0] p48_add_68510_comb;
  wire [31:0] p48_add_68512_comb;
  wire [31:0] p48_add_68530_comb;
  wire [31:0] p48_add_68513_comb;
  wire [31:0] p48_add_68531_comb;
  assign p48_add_68510_comb = {p47_add_68398[5:0] ^ p47_add_68398[10:5] ^ p47_add_68398[24:19], p47_add_68398[31:27] ^ p47_add_68398[4:0] ^ p47_add_68398[18:14], p47_add_68398[26:13] ^ p47_add_68398[31:18] ^ p47_add_68398[13:0], p47_add_68398[12:6] ^ p47_add_68398[17:11] ^ p47_add_68398[31:25]} + (p47_add_68398 & p47_add_68262 ^ ~(p47_add_68398 | ~p47_add_68109));
  assign p48_add_68512_comb = p48_add_68510_comb + 32'ha81a_664b;
  assign p48_add_68530_comb = p47_add_67524 + {p47_add_68438[16:7] ^ p47_add_68438[18:9], p47_add_68438[6:0] ^ p47_add_68438[8:2] ^ p47_add_68438[31:25], p47_add_68438[31:30] ^ p47_add_68438[1:0] ^ p47_add_68438[24:23], p47_add_68438[29:17] ^ p47_add_68438[31:19] ^ p47_add_68438[22:10]};
  assign p48_add_68513_comb = p48_add_68512_comb + p47_add_68285;
  assign p48_add_68531_comb = p47_add_67903 + p48_add_68530_comb;

  // Registers for pipe stage 48:
  reg [31:0] p48_add_68109;
  reg [31:0] p48_add_68262;
  reg [31:0] p48_add_68398;
  reg [31:0] p48_add_68022;
  reg [31:0] p48_add_68513;
  reg [31:0] p48_add_68156;
  reg [31:0] p48_add_68307;
  reg [31:0] p48_and_68415;
  reg [31:0] p48_add_68420;
  reg [31:0] p48_add_68342;
  reg [31:0] p48_add_68208;
  reg [31:0] p48_add_68191;
  reg [31:0] p48_add_68058;
  reg [31:0] p48_add_68041;
  reg [31:0] p48_add_68531;
  reg [31:0] p48_add_67886;
  reg [31:0] p48_add_68438;
  reg [31:0] p48_add_67741;
  reg [31:0] p48_add_68325;
  reg [31:0] p48_add_67869;
  reg [31:0] p48_add_68174;
  reg [31:0] p48_add_67524;
  reg [31:0] p48_add_68024;
  reg [31:0] p48_add_66624;
  reg [31:0] p48_add_67851;
  always_ff @ (posedge clk) begin
    p48_add_68109 <= p47_add_68109;
    p48_add_68262 <= p47_add_68262;
    p48_add_68398 <= p47_add_68398;
    p48_add_68022 <= p47_add_68022;
    p48_add_68513 <= p48_add_68513_comb;
    p48_add_68156 <= p47_add_68156;
    p48_add_68307 <= p47_add_68307;
    p48_and_68415 <= p47_and_68415;
    p48_add_68420 <= p47_add_68420;
    p48_add_68342 <= p47_add_68342;
    p48_add_68208 <= p47_add_68208;
    p48_add_68191 <= p47_add_68191;
    p48_add_68058 <= p47_add_68058;
    p48_add_68041 <= p47_add_68041;
    p48_add_68531 <= p48_add_68531_comb;
    p48_add_67886 <= p47_add_67886;
    p48_add_68438 <= p47_add_68438;
    p48_add_67741 <= p47_add_67741;
    p48_add_68325 <= p47_add_68325;
    p48_add_67869 <= p47_add_67869;
    p48_add_68174 <= p47_add_68174;
    p48_add_67524 <= p47_add_67524;
    p48_add_68024 <= p47_add_68024;
    p48_add_66624 <= p47_add_66624;
    p48_add_67851 <= p47_add_67851;
  end

  // ===== Pipe stage 49:
  wire [31:0] p49_add_68582_comb;
  wire [1:0] p49_bit_slice_68631_comb;
  wire [31:0] p49_and_68629_comb;
  wire [27:0] p49_add_68604_comb;
  wire [31:0] p49_add_68634_comb;
  wire [31:0] p49_add_68651_comb;
  wire [31:0] p49_add_68609_comb;
  wire [31:0] p49_add_68610_comb;
  wire [31:0] p49_add_68612_comb;
  wire [31:0] p49_add_68635_comb;
  wire [31:0] p49_add_68685_comb;
  wire [31:0] p49_add_68669_comb;
  wire [31:0] p49_add_68652_comb;
  wire [31:0] p49_add_68611_comb;
  assign p49_add_68582_comb = p48_add_68022 + p48_add_68513;
  assign p49_bit_slice_68631_comb = p48_add_67869[1:0];
  assign p49_and_68629_comb = p48_add_68420 & p48_add_68307;
  assign p49_add_68604_comb = p48_add_68024[31:4] + 28'hc24_b8b7;
  assign p49_add_68634_comb = {p48_add_68420[1:0] ^ p48_add_68420[12:11] ^ p48_add_68420[21:20], p48_add_68420[31:21] ^ p48_add_68420[10:0] ^ p48_add_68420[19:9], p48_add_68420[20:12] ^ p48_add_68420[31:23] ^ p48_add_68420[8:0], p48_add_68420[11:2] ^ p48_add_68420[22:13] ^ p48_add_68420[31:22]} + (p49_and_68629_comb ^ p48_add_68420 & p48_add_68156 ^ p48_and_68415);
  assign p49_add_68651_comb = p48_add_67851 + {p48_add_67869[16:7] ^ p48_add_67869[18:9], p48_add_67869[6:0] ^ p48_add_67869[8:2] ^ p48_add_67869[31:25], p48_add_67869[31:30] ^ p49_bit_slice_68631_comb ^ p48_add_67869[24:23], p48_add_67869[29:17] ^ p48_add_67869[31:19] ^ p48_add_67869[22:10]};
  assign p49_add_68609_comb = {p49_add_68582_comb[5:0] ^ p49_add_68582_comb[10:5] ^ p49_add_68582_comb[24:19], p49_add_68582_comb[31:27] ^ p49_add_68582_comb[4:0] ^ p49_add_68582_comb[18:14], p49_add_68582_comb[26:13] ^ p49_add_68582_comb[31:18] ^ p49_add_68582_comb[13:0], p49_add_68582_comb[12:6] ^ p49_add_68582_comb[17:11] ^ p49_add_68582_comb[31:25]} + p48_add_68109;
  assign p49_add_68610_comb = (p49_add_68582_comb & p48_add_68398 ^ ~(p49_add_68582_comb | ~p48_add_68262)) + {p49_add_68604_comb, p48_add_68024[3:0]};
  assign p49_add_68612_comb = p48_add_68262 + p48_add_67524;
  assign p49_add_68635_comb = p48_add_68513 + p49_add_68634_comb;
  assign p49_add_68685_comb = {p48_add_68024[6:4] ^ p48_add_68024[17:15], p48_add_68024[3:0] ^ p48_add_68024[14:11] ^ p48_add_68024[31:28], p48_add_68024[31:21] ^ p48_add_68024[10:0] ^ p48_add_68024[27:17], p48_add_68024[20:7] ^ p48_add_68024[31:18] ^ p48_add_68024[16:3]} + p48_add_66624;
  assign p49_add_68669_comb = {p48_add_66624[6:4] ^ p48_add_66624[17:15], p48_add_66624[3:0] ^ p48_add_66624[14:11] ^ p48_add_66624[31:28], p48_add_66624[31:21] ^ p48_add_66624[10:0] ^ p48_add_66624[27:17], p48_add_66624[20:7] ^ p48_add_66624[31:18] ^ p48_add_66624[16:3]} + p48_add_67851;
  assign p49_add_68652_comb = p48_add_67741 + p49_add_68651_comb;
  assign p49_add_68611_comb = p49_add_68609_comb + p49_add_68610_comb;

  // Registers for pipe stage 49:
  reg [31:0] p49_add_68398;
  reg [31:0] p49_add_68582;
  reg [31:0] p49_add_68156;
  reg [31:0] p49_add_68612;
  reg [31:0] p49_add_68307;
  reg [31:0] p49_add_68420;
  reg [1:0] p49_bit_slice_68631;
  reg [31:0] p49_and_68629;
  reg [31:0] p49_add_68635;
  reg [31:0] p49_add_68685;
  reg [31:0] p49_add_68669;
  reg [31:0] p49_add_68342;
  reg [31:0] p49_add_68208;
  reg [31:0] p49_add_68191;
  reg [31:0] p49_add_68058;
  reg [31:0] p49_add_68041;
  reg [31:0] p49_add_68531;
  reg [31:0] p49_add_67886;
  reg [31:0] p49_add_68438;
  reg [31:0] p49_add_68652;
  reg [31:0] p49_add_68325;
  reg [31:0] p49_add_67869;
  reg [31:0] p49_add_68174;
  reg [31:0] p49_add_67524;
  reg [31:0] p49_add_68611;
  reg [31:0] p49_add_68024;
  always_ff @ (posedge clk) begin
    p49_add_68398 <= p48_add_68398;
    p49_add_68582 <= p49_add_68582_comb;
    p49_add_68156 <= p48_add_68156;
    p49_add_68612 <= p49_add_68612_comb;
    p49_add_68307 <= p48_add_68307;
    p49_add_68420 <= p48_add_68420;
    p49_bit_slice_68631 <= p49_bit_slice_68631_comb;
    p49_and_68629 <= p49_and_68629_comb;
    p49_add_68635 <= p49_add_68635_comb;
    p49_add_68685 <= p49_add_68685_comb;
    p49_add_68669 <= p49_add_68669_comb;
    p49_add_68342 <= p48_add_68342;
    p49_add_68208 <= p48_add_68208;
    p49_add_68191 <= p48_add_68191;
    p49_add_68058 <= p48_add_68058;
    p49_add_68041 <= p48_add_68041;
    p49_add_68531 <= p48_add_68531;
    p49_add_67886 <= p48_add_67886;
    p49_add_68438 <= p48_add_68438;
    p49_add_68652 <= p49_add_68652_comb;
    p49_add_68325 <= p48_add_68325;
    p49_add_67869 <= p48_add_67869;
    p49_add_68174 <= p48_add_68174;
    p49_add_67524 <= p48_add_67524;
    p49_add_68611 <= p49_add_68611_comb;
    p49_add_68024 <= p48_add_68024;
  end

  // ===== Pipe stage 50:
  wire [31:0] p50_add_68738_comb;
  wire [31:0] p50_and_68780_comb;
  wire [31:0] p50_add_68784_comb;
  wire [31:0] p50_add_68760_comb;
  wire [31:0] p50_add_68802_comb;
  wire [31:0] p50_add_68763_comb;
  wire [31:0] p50_add_68785_comb;
  wire [31:0] p50_add_68762_comb;
  wire [31:0] p50_add_68837_comb;
  wire [31:0] p50_add_68820_comb;
  wire [31:0] p50_add_68803_comb;
  assign p50_add_68738_comb = p49_add_68156 + p49_add_68611;
  assign p50_and_68780_comb = p49_add_68635 & p49_add_68420;
  assign p50_add_68784_comb = {p49_add_68635[1:0] ^ p49_add_68635[12:11] ^ p49_add_68635[21:20], p49_add_68635[31:21] ^ p49_add_68635[10:0] ^ p49_add_68635[19:9], p49_add_68635[20:12] ^ p49_add_68635[31:23] ^ p49_add_68635[8:0], p49_add_68635[11:2] ^ p49_add_68635[22:13] ^ p49_add_68635[31:22]} + (p50_and_68780_comb ^ p49_add_68635 & p49_add_68307 ^ p49_and_68629);
  assign p50_add_68760_comb = {p50_add_68738_comb[5:0] ^ p50_add_68738_comb[10:5] ^ p50_add_68738_comb[24:19], p50_add_68738_comb[31:27] ^ p50_add_68738_comb[4:0] ^ p50_add_68738_comb[18:14], p50_add_68738_comb[26:13] ^ p50_add_68738_comb[31:18] ^ p50_add_68738_comb[13:0], p50_add_68738_comb[12:6] ^ p50_add_68738_comb[17:11] ^ p50_add_68738_comb[31:25]} + (p50_add_68738_comb & p49_add_68582 ^ ~(p50_add_68738_comb | ~p49_add_68398));
  assign p50_add_68802_comb = p49_add_68024 + {p49_add_68652[16:7] ^ p49_add_68652[18:9], p49_add_68652[6:0] ^ p49_add_68652[8:2] ^ p49_add_68652[31:25], p49_add_68652[31:30] ^ p49_add_68652[1:0] ^ p49_add_68652[24:23], p49_add_68652[29:17] ^ p49_add_68652[31:19] ^ p49_add_68652[22:10]};
  assign p50_add_68763_comb = p49_add_68398 + p49_add_68174;
  assign p50_add_68785_comb = p49_add_68611 + p50_add_68784_comb;
  assign p50_add_68762_comb = p50_add_68760_comb + 32'hc76c_51a3;
  assign p50_add_68837_comb = {p49_add_68174[6:4] ^ p49_add_68174[17:15], p49_add_68174[3:0] ^ p49_add_68174[14:11] ^ p49_add_68174[31:28], p49_add_68174[31:21] ^ p49_add_68174[10:0] ^ p49_add_68174[27:17], p49_add_68174[20:7] ^ p49_add_68174[31:18] ^ p49_add_68174[16:3]} + p49_add_67524;
  assign p50_add_68820_comb = {p49_add_67524[6:4] ^ p49_add_67524[17:15], p49_add_67524[3:0] ^ p49_add_67524[14:11] ^ p49_add_67524[31:28], p49_add_67524[31:21] ^ p49_add_67524[10:0] ^ p49_add_67524[27:17], p49_add_67524[20:7] ^ p49_add_67524[31:18] ^ p49_add_67524[16:3]} + p49_add_68024;
  assign p50_add_68803_comb = p49_add_67886 + p50_add_68802_comb;

  // Registers for pipe stage 50:
  reg [31:0] p50_add_68582;
  reg [31:0] p50_add_68738;
  reg [31:0] p50_add_68612;
  reg [31:0] p50_add_68307;
  reg [31:0] p50_add_68763;
  reg [31:0] p50_add_68420;
  reg [1:0] p50_bit_slice_68631;
  reg [31:0] p50_add_68635;
  reg [31:0] p50_and_68780;
  reg [31:0] p50_add_68785;
  reg [31:0] p50_add_68762;
  reg [31:0] p50_add_68837;
  reg [31:0] p50_add_68820;
  reg [31:0] p50_add_68685;
  reg [31:0] p50_add_68669;
  reg [31:0] p50_add_68342;
  reg [31:0] p50_add_68208;
  reg [31:0] p50_add_68191;
  reg [31:0] p50_add_68058;
  reg [31:0] p50_add_68041;
  reg [31:0] p50_add_68531;
  reg [31:0] p50_add_68803;
  reg [31:0] p50_add_68438;
  reg [31:0] p50_add_68652;
  reg [31:0] p50_add_68325;
  reg [31:0] p50_add_67869;
  reg [31:0] p50_add_68174;
  always_ff @ (posedge clk) begin
    p50_add_68582 <= p49_add_68582;
    p50_add_68738 <= p50_add_68738_comb;
    p50_add_68612 <= p49_add_68612;
    p50_add_68307 <= p49_add_68307;
    p50_add_68763 <= p50_add_68763_comb;
    p50_add_68420 <= p49_add_68420;
    p50_bit_slice_68631 <= p49_bit_slice_68631;
    p50_add_68635 <= p49_add_68635;
    p50_and_68780 <= p50_and_68780_comb;
    p50_add_68785 <= p50_add_68785_comb;
    p50_add_68762 <= p50_add_68762_comb;
    p50_add_68837 <= p50_add_68837_comb;
    p50_add_68820 <= p50_add_68820_comb;
    p50_add_68685 <= p49_add_68685;
    p50_add_68669 <= p49_add_68669;
    p50_add_68342 <= p49_add_68342;
    p50_add_68208 <= p49_add_68208;
    p50_add_68191 <= p49_add_68191;
    p50_add_68058 <= p49_add_68058;
    p50_add_68041 <= p49_add_68041;
    p50_add_68531 <= p49_add_68531;
    p50_add_68803 <= p50_add_68803_comb;
    p50_add_68438 <= p49_add_68438;
    p50_add_68652 <= p49_add_68652;
    p50_add_68325 <= p49_add_68325;
    p50_add_67869 <= p49_add_67869;
    p50_add_68174 <= p49_add_68174;
  end

  // ===== Pipe stage 51:
  wire [31:0] p51_add_68892_comb;
  wire [31:0] p51_add_68893_comb;
  wire [31:0] p51_and_68932_comb;
  wire [31:0] p51_add_68936_comb;
  wire [31:0] p51_add_68954_comb;
  wire [31:0] p51_add_68915_comb;
  wire [31:0] p51_add_68937_comb;
  wire [31:0] p51_add_68972_comb;
  wire [31:0] p51_add_68955_comb;
  assign p51_add_68892_comb = p50_add_68762 + p50_add_68612;
  assign p51_add_68893_comb = p50_add_68307 + p51_add_68892_comb;
  assign p51_and_68932_comb = p50_add_68785 & p50_add_68635;
  assign p51_add_68936_comb = {p50_add_68785[1:0] ^ p50_add_68785[12:11] ^ p50_add_68785[21:20], p50_add_68785[31:21] ^ p50_add_68785[10:0] ^ p50_add_68785[19:9], p50_add_68785[20:12] ^ p50_add_68785[31:23] ^ p50_add_68785[8:0], p50_add_68785[11:2] ^ p50_add_68785[22:13] ^ p50_add_68785[31:22]} + (p51_and_68932_comb ^ p50_add_68785 & p50_add_68420 ^ p50_and_68780);
  assign p51_add_68954_comb = p50_add_68174 + {p50_add_68803[16:7] ^ p50_add_68803[18:9], p50_add_68803[6:0] ^ p50_add_68803[8:2] ^ p50_add_68803[31:25], p50_add_68803[31:30] ^ p50_add_68803[1:0] ^ p50_add_68803[24:23], p50_add_68803[29:17] ^ p50_add_68803[31:19] ^ p50_add_68803[22:10]};
  assign p51_add_68915_comb = {p51_add_68893_comb[5:0] ^ p51_add_68893_comb[10:5] ^ p51_add_68893_comb[24:19], p51_add_68893_comb[31:27] ^ p51_add_68893_comb[4:0] ^ p51_add_68893_comb[18:14], p51_add_68893_comb[26:13] ^ p51_add_68893_comb[31:18] ^ p51_add_68893_comb[13:0], p51_add_68893_comb[12:6] ^ p51_add_68893_comb[17:11] ^ p51_add_68893_comb[31:25]} + (p51_add_68893_comb & p50_add_68738 ^ ~(p51_add_68893_comb | ~p50_add_68582));
  assign p51_add_68937_comb = p51_add_68892_comb + p51_add_68936_comb;
  assign p51_add_68972_comb = {p50_add_67869[6:4] ^ p50_add_67869[17:15], p50_add_67869[3:0] ^ p50_add_67869[14:11] ^ p50_add_67869[31:28], p50_add_67869[31:21] ^ p50_add_67869[10:0] ^ p50_add_67869[27:17], p50_add_67869[20:7] ^ p50_add_67869[31:18] ^ p50_add_67869[16:3]} + p50_add_68174;
  assign p51_add_68955_comb = p50_add_68041 + p51_add_68954_comb;

  // Registers for pipe stage 51:
  reg [31:0] p51_add_68582;
  reg [31:0] p51_add_68738;
  reg [31:0] p51_add_68893;
  reg [31:0] p51_add_68915;
  reg [31:0] p51_add_68763;
  reg [31:0] p51_add_68420;
  reg [1:0] p51_bit_slice_68631;
  reg [31:0] p51_add_68635;
  reg [31:0] p51_add_68785;
  reg [31:0] p51_and_68932;
  reg [31:0] p51_add_68937;
  reg [31:0] p51_add_68972;
  reg [31:0] p51_add_68837;
  reg [31:0] p51_add_68820;
  reg [31:0] p51_add_68685;
  reg [31:0] p51_add_68669;
  reg [31:0] p51_add_68342;
  reg [31:0] p51_add_68208;
  reg [31:0] p51_add_68191;
  reg [31:0] p51_add_68058;
  reg [31:0] p51_add_68955;
  reg [31:0] p51_add_68531;
  reg [31:0] p51_add_68803;
  reg [31:0] p51_add_68438;
  reg [31:0] p51_add_68652;
  reg [31:0] p51_add_68325;
  reg [31:0] p51_add_67869;
  always_ff @ (posedge clk) begin
    p51_add_68582 <= p50_add_68582;
    p51_add_68738 <= p50_add_68738;
    p51_add_68893 <= p51_add_68893_comb;
    p51_add_68915 <= p51_add_68915_comb;
    p51_add_68763 <= p50_add_68763;
    p51_add_68420 <= p50_add_68420;
    p51_bit_slice_68631 <= p50_bit_slice_68631;
    p51_add_68635 <= p50_add_68635;
    p51_add_68785 <= p50_add_68785;
    p51_and_68932 <= p51_and_68932_comb;
    p51_add_68937 <= p51_add_68937_comb;
    p51_add_68972 <= p51_add_68972_comb;
    p51_add_68837 <= p50_add_68837;
    p51_add_68820 <= p50_add_68820;
    p51_add_68685 <= p50_add_68685;
    p51_add_68669 <= p50_add_68669;
    p51_add_68342 <= p50_add_68342;
    p51_add_68208 <= p50_add_68208;
    p51_add_68191 <= p50_add_68191;
    p51_add_68058 <= p50_add_68058;
    p51_add_68955 <= p51_add_68955_comb;
    p51_add_68531 <= p50_add_68531;
    p51_add_68803 <= p50_add_68803;
    p51_add_68438 <= p50_add_68438;
    p51_add_68652 <= p50_add_68652;
    p51_add_68325 <= p50_add_68325;
    p51_add_67869 <= p50_add_67869;
  end

  // ===== Pipe stage 52:
  wire [31:0] p52_and_69051_comb;
  wire [31:0] p52_add_69028_comb;
  wire [31:0] p52_add_69029_comb;
  wire [29:0] p52_add_69033_comb;
  wire [31:0] p52_add_69055_comb;
  wire [31:0] p52_add_69073_comb;
  wire [31:0] p52_add_69030_comb;
  wire [31:0] p52_concat_69034_comb;
  wire [31:0] p52_add_69056_comb;
  wire [31:0] p52_add_69074_comb;
  assign p52_and_69051_comb = p51_add_68937 & p51_add_68785;
  assign p52_add_69028_comb = p51_add_68915 + 32'hd192_e819;
  assign p52_add_69029_comb = p52_add_69028_comb + p51_add_68763;
  assign p52_add_69033_comb = p51_add_67869[31:2] + 30'h35a6_4189;
  assign p52_add_69055_comb = {p51_add_68937[1:0] ^ p51_add_68937[12:11] ^ p51_add_68937[21:20], p51_add_68937[31:21] ^ p51_add_68937[10:0] ^ p51_add_68937[19:9], p51_add_68937[20:12] ^ p51_add_68937[31:23] ^ p51_add_68937[8:0], p51_add_68937[11:2] ^ p51_add_68937[22:13] ^ p51_add_68937[31:22]} + (p52_and_69051_comb ^ p51_add_68937 & p51_add_68635 ^ p51_and_68932);
  assign p52_add_69073_comb = p51_add_68325 + {p51_add_68955[16:7] ^ p51_add_68955[18:9], p51_add_68955[6:0] ^ p51_add_68955[8:2] ^ p51_add_68955[31:25], p51_add_68955[31:30] ^ p51_add_68955[1:0] ^ p51_add_68955[24:23], p51_add_68955[29:17] ^ p51_add_68955[31:19] ^ p51_add_68955[22:10]};
  assign p52_add_69030_comb = p51_add_68420 + p52_add_69029_comb;
  assign p52_concat_69034_comb = {p52_add_69033_comb, p51_bit_slice_68631};
  assign p52_add_69056_comb = p52_add_69029_comb + p52_add_69055_comb;
  assign p52_add_69074_comb = p51_add_68191 + p52_add_69073_comb;

  // Registers for pipe stage 52:
  reg [31:0] p52_add_68582;
  reg [31:0] p52_add_68738;
  reg [31:0] p52_add_68893;
  reg [31:0] p52_add_69030;
  reg [31:0] p52_concat_69034;
  reg [31:0] p52_add_68635;
  reg [31:0] p52_add_68785;
  reg [31:0] p52_add_68937;
  reg [31:0] p52_and_69051;
  reg [31:0] p52_add_69056;
  reg [31:0] p52_add_68972;
  reg [31:0] p52_add_68837;
  reg [31:0] p52_add_68820;
  reg [31:0] p52_add_68685;
  reg [31:0] p52_add_68669;
  reg [31:0] p52_add_68342;
  reg [31:0] p52_add_68208;
  reg [31:0] p52_add_69074;
  reg [31:0] p52_add_68058;
  reg [31:0] p52_add_68955;
  reg [31:0] p52_add_68531;
  reg [31:0] p52_add_68803;
  reg [31:0] p52_add_68438;
  reg [31:0] p52_add_68652;
  reg [31:0] p52_add_68325;
  reg [31:0] p52_add_67869;
  always_ff @ (posedge clk) begin
    p52_add_68582 <= p51_add_68582;
    p52_add_68738 <= p51_add_68738;
    p52_add_68893 <= p51_add_68893;
    p52_add_69030 <= p52_add_69030_comb;
    p52_concat_69034 <= p52_concat_69034_comb;
    p52_add_68635 <= p51_add_68635;
    p52_add_68785 <= p51_add_68785;
    p52_add_68937 <= p51_add_68937;
    p52_and_69051 <= p52_and_69051_comb;
    p52_add_69056 <= p52_add_69056_comb;
    p52_add_68972 <= p51_add_68972;
    p52_add_68837 <= p51_add_68837;
    p52_add_68820 <= p51_add_68820;
    p52_add_68685 <= p51_add_68685;
    p52_add_68669 <= p51_add_68669;
    p52_add_68342 <= p51_add_68342;
    p52_add_68208 <= p51_add_68208;
    p52_add_69074 <= p52_add_69074_comb;
    p52_add_68058 <= p51_add_68058;
    p52_add_68955 <= p51_add_68955;
    p52_add_68531 <= p51_add_68531;
    p52_add_68803 <= p51_add_68803;
    p52_add_68438 <= p51_add_68438;
    p52_add_68652 <= p51_add_68652;
    p52_add_68325 <= p51_add_68325;
    p52_add_67869 <= p51_add_67869;
  end

  // ===== Pipe stage 53:
  wire [31:0] p53_and_69169_comb;
  wire [31:0] p53_add_69148_comb;
  wire [31:0] p53_add_69149_comb;
  wire [31:0] p53_add_69150_comb;
  wire [31:0] p53_add_69173_comb;
  wire [31:0] p53_add_69191_comb;
  wire [31:0] p53_add_69151_comb;
  wire [31:0] p53_add_69152_comb;
  wire [31:0] p53_add_69174_comb;
  wire [31:0] p53_add_69192_comb;
  assign p53_and_69169_comb = p52_add_69056 & p52_add_68937;
  assign p53_add_69148_comb = {p52_add_69030[5:0] ^ p52_add_69030[10:5] ^ p52_add_69030[24:19], p52_add_69030[31:27] ^ p52_add_69030[4:0] ^ p52_add_69030[18:14], p52_add_69030[26:13] ^ p52_add_69030[31:18] ^ p52_add_69030[13:0], p52_add_69030[12:6] ^ p52_add_69030[17:11] ^ p52_add_69030[31:25]} + p52_add_68582;
  assign p53_add_69149_comb = (p52_add_69030 & p52_add_68893 ^ ~(p52_add_69030 | ~p52_add_68738)) + p52_concat_69034;
  assign p53_add_69150_comb = p53_add_69148_comb + p53_add_69149_comb;
  assign p53_add_69173_comb = {p52_add_69056[1:0] ^ p52_add_69056[12:11] ^ p52_add_69056[21:20], p52_add_69056[31:21] ^ p52_add_69056[10:0] ^ p52_add_69056[19:9], p52_add_69056[20:12] ^ p52_add_69056[31:23] ^ p52_add_69056[8:0], p52_add_69056[11:2] ^ p52_add_69056[22:13] ^ p52_add_69056[31:22]} + (p53_and_69169_comb ^ p52_add_69056 & p52_add_68785 ^ p52_and_69051);
  assign p53_add_69191_comb = p52_add_68438 + {p52_add_69074[16:7] ^ p52_add_69074[18:9], p52_add_69074[6:0] ^ p52_add_69074[8:2] ^ p52_add_69074[31:25], p52_add_69074[31:30] ^ p52_add_69074[1:0] ^ p52_add_69074[24:23], p52_add_69074[29:17] ^ p52_add_69074[31:19] ^ p52_add_69074[22:10]};
  assign p53_add_69151_comb = p52_add_68635 + p53_add_69150_comb;
  assign p53_add_69152_comb = p52_add_68738 + p52_add_68325;
  assign p53_add_69174_comb = p53_add_69150_comb + p53_add_69173_comb;
  assign p53_add_69192_comb = p52_add_68342 + p53_add_69191_comb;

  // Registers for pipe stage 53:
  reg [31:0] p53_add_68893;
  reg [31:0] p53_add_69030;
  reg [31:0] p53_add_69151;
  reg [31:0] p53_add_69152;
  reg [31:0] p53_add_68785;
  reg [31:0] p53_add_68937;
  reg [31:0] p53_add_69056;
  reg [31:0] p53_and_69169;
  reg [31:0] p53_add_69174;
  reg [31:0] p53_add_68972;
  reg [31:0] p53_add_68837;
  reg [31:0] p53_add_68820;
  reg [31:0] p53_add_68685;
  reg [31:0] p53_add_68669;
  reg [31:0] p53_add_69192;
  reg [31:0] p53_add_68208;
  reg [31:0] p53_add_69074;
  reg [31:0] p53_add_68058;
  reg [31:0] p53_add_68955;
  reg [31:0] p53_add_68531;
  reg [31:0] p53_add_68803;
  reg [31:0] p53_add_68438;
  reg [31:0] p53_add_68652;
  reg [31:0] p53_add_68325;
  reg [31:0] p53_add_67869;
  always_ff @ (posedge clk) begin
    p53_add_68893 <= p52_add_68893;
    p53_add_69030 <= p52_add_69030;
    p53_add_69151 <= p53_add_69151_comb;
    p53_add_69152 <= p53_add_69152_comb;
    p53_add_68785 <= p52_add_68785;
    p53_add_68937 <= p52_add_68937;
    p53_add_69056 <= p52_add_69056;
    p53_and_69169 <= p53_and_69169_comb;
    p53_add_69174 <= p53_add_69174_comb;
    p53_add_68972 <= p52_add_68972;
    p53_add_68837 <= p52_add_68837;
    p53_add_68820 <= p52_add_68820;
    p53_add_68685 <= p52_add_68685;
    p53_add_68669 <= p52_add_68669;
    p53_add_69192 <= p53_add_69192_comb;
    p53_add_68208 <= p52_add_68208;
    p53_add_69074 <= p52_add_69074;
    p53_add_68058 <= p52_add_68058;
    p53_add_68955 <= p52_add_68955;
    p53_add_68531 <= p52_add_68531;
    p53_add_68803 <= p52_add_68803;
    p53_add_68438 <= p52_add_68438;
    p53_add_68652 <= p52_add_68652;
    p53_add_68325 <= p52_add_68325;
    p53_add_67869 <= p52_add_67869;
  end

  // ===== Pipe stage 54:
  wire [31:0] p54_add_69264_comb;
  wire [31:0] p54_add_69266_comb;
  wire [29:0] p54_add_69270_comb;
  wire [31:0] p54_add_69306_comb;
  wire [31:0] p54_add_69288_comb;
  wire [31:0] p54_add_69267_comb;
  wire [31:0] p54_concat_69272_comb;
  wire [31:0] p54_add_69324_comb;
  wire [31:0] p54_add_69307_comb;
  wire [31:0] p54_add_69289_comb;
  assign p54_add_69264_comb = {p53_add_69151[5:0] ^ p53_add_69151[10:5] ^ p53_add_69151[24:19], p53_add_69151[31:27] ^ p53_add_69151[4:0] ^ p53_add_69151[18:14], p53_add_69151[26:13] ^ p53_add_69151[31:18] ^ p53_add_69151[13:0], p53_add_69151[12:6] ^ p53_add_69151[17:11] ^ p53_add_69151[31:25]} + (p53_add_69151 & p53_add_69030 ^ ~(p53_add_69151 | ~p53_add_68893));
  assign p54_add_69266_comb = p54_add_69264_comb + 32'hf40e_3585;
  assign p54_add_69270_comb = p53_add_68531[31:2] + 30'h09d2_1dd3;
  assign p54_add_69306_comb = p53_add_68531 + {p53_add_69192[16:7] ^ p53_add_69192[18:9], p53_add_69192[6:0] ^ p53_add_69192[8:2] ^ p53_add_69192[31:25], p53_add_69192[31:30] ^ p53_add_69192[1:0] ^ p53_add_69192[24:23], p53_add_69192[29:17] ^ p53_add_69192[31:19] ^ p53_add_69192[22:10]};
  assign p54_add_69288_comb = p53_add_67869 + {p53_add_68531[16:7] ^ p53_add_68531[18:9], p53_add_68531[6:0] ^ p53_add_68531[8:2] ^ p53_add_68531[31:25], p53_add_68531[31:30] ^ p53_add_68531[1:0] ^ p53_add_68531[24:23], p53_add_68531[29:17] ^ p53_add_68531[31:19] ^ p53_add_68531[22:10]};
  assign p54_add_69267_comb = p54_add_69266_comb + p53_add_69152;
  assign p54_concat_69272_comb = {p54_add_69270_comb, p53_add_68531[1:0]};
  assign p54_add_69324_comb = {p53_add_68325[6:4] ^ p53_add_68325[17:15], p53_add_68325[3:0] ^ p53_add_68325[14:11] ^ p53_add_68325[31:28], p53_add_68325[31:21] ^ p53_add_68325[10:0] ^ p53_add_68325[27:17], p53_add_68325[20:7] ^ p53_add_68325[31:18] ^ p53_add_68325[16:3]} + p53_add_67869;
  assign p54_add_69307_comb = p53_add_68685 + p54_add_69306_comb;
  assign p54_add_69289_comb = p53_add_68058 + p54_add_69288_comb;

  // Registers for pipe stage 54:
  reg [31:0] p54_add_68893;
  reg [31:0] p54_add_69030;
  reg [31:0] p54_add_69151;
  reg [31:0] p54_add_68785;
  reg [31:0] p54_add_69267;
  reg [31:0] p54_add_68937;
  reg [31:0] p54_add_69056;
  reg [31:0] p54_and_69169;
  reg [31:0] p54_add_69174;
  reg [31:0] p54_concat_69272;
  reg [31:0] p54_add_69324;
  reg [31:0] p54_add_68972;
  reg [31:0] p54_add_68837;
  reg [31:0] p54_add_68820;
  reg [31:0] p54_add_69307;
  reg [31:0] p54_add_68669;
  reg [31:0] p54_add_69192;
  reg [31:0] p54_add_68208;
  reg [31:0] p54_add_69074;
  reg [31:0] p54_add_69289;
  reg [31:0] p54_add_68955;
  reg [31:0] p54_add_68803;
  reg [31:0] p54_add_68438;
  reg [31:0] p54_add_68652;
  reg [31:0] p54_add_68325;
  always_ff @ (posedge clk) begin
    p54_add_68893 <= p53_add_68893;
    p54_add_69030 <= p53_add_69030;
    p54_add_69151 <= p53_add_69151;
    p54_add_68785 <= p53_add_68785;
    p54_add_69267 <= p54_add_69267_comb;
    p54_add_68937 <= p53_add_68937;
    p54_add_69056 <= p53_add_69056;
    p54_and_69169 <= p53_and_69169;
    p54_add_69174 <= p53_add_69174;
    p54_concat_69272 <= p54_concat_69272_comb;
    p54_add_69324 <= p54_add_69324_comb;
    p54_add_68972 <= p53_add_68972;
    p54_add_68837 <= p53_add_68837;
    p54_add_68820 <= p53_add_68820;
    p54_add_69307 <= p54_add_69307_comb;
    p54_add_68669 <= p53_add_68669;
    p54_add_69192 <= p53_add_69192;
    p54_add_68208 <= p53_add_68208;
    p54_add_69074 <= p53_add_69074;
    p54_add_69289 <= p54_add_69289_comb;
    p54_add_68955 <= p53_add_68955;
    p54_add_68803 <= p53_add_68803;
    p54_add_68438 <= p53_add_68438;
    p54_add_68652 <= p53_add_68652;
    p54_add_68325 <= p53_add_68325;
  end

  // ===== Pipe stage 55:
  wire [31:0] p55_add_69375_comb;
  wire [31:0] p55_and_69421_comb;
  wire [27:0] p55_add_69397_comb;
  wire [31:0] p55_add_69425_comb;
  wire [31:0] p55_add_69461_comb;
  wire [31:0] p55_add_69443_comb;
  wire [31:0] p55_add_69402_comb;
  wire [31:0] p55_add_69403_comb;
  wire [31:0] p55_add_69426_comb;
  wire [3:0] p55_xor_69465_comb;
  wire [31:0] p55_add_69462_comb;
  wire [31:0] p55_add_69444_comb;
  wire [31:0] p55_add_69404_comb;
  assign p55_add_69375_comb = p54_add_68785 + p54_add_69267;
  assign p55_and_69421_comb = p54_add_69174 & p54_add_69056;
  assign p55_add_69397_comb = p54_add_68652[31:4] + 28'h106_aa07;
  assign p55_add_69425_comb = {p54_add_69174[1:0] ^ p54_add_69174[12:11] ^ p54_add_69174[21:20], p54_add_69174[31:21] ^ p54_add_69174[10:0] ^ p54_add_69174[19:9], p54_add_69174[20:12] ^ p54_add_69174[31:23] ^ p54_add_69174[8:0], p54_add_69174[11:2] ^ p54_add_69174[22:13] ^ p54_add_69174[31:22]} + (p55_and_69421_comb ^ p54_add_69174 & p54_add_68937 ^ p54_and_69169);
  assign p55_add_69461_comb = p54_add_69289 + {p54_add_69307[16:7] ^ p54_add_69307[18:9], p54_add_69307[6:0] ^ p54_add_69307[8:2] ^ p54_add_69307[31:25], p54_add_69307[31:30] ^ p54_add_69307[1:0] ^ p54_add_69307[24:23], p54_add_69307[29:17] ^ p54_add_69307[31:19] ^ p54_add_69307[22:10]};
  assign p55_add_69443_comb = p54_add_68652 + {p54_add_69289[16:7] ^ p54_add_69289[18:9], p54_add_69289[6:0] ^ p54_add_69289[8:2] ^ p54_add_69289[31:25], p54_add_69289[31:30] ^ p54_add_69289[1:0] ^ p54_add_69289[24:23], p54_add_69289[29:17] ^ p54_add_69289[31:19] ^ p54_add_69289[22:10]};
  assign p55_add_69402_comb = {p55_add_69375_comb[5:0] ^ p55_add_69375_comb[10:5] ^ p55_add_69375_comb[24:19], p55_add_69375_comb[31:27] ^ p55_add_69375_comb[4:0] ^ p55_add_69375_comb[18:14], p55_add_69375_comb[26:13] ^ p55_add_69375_comb[31:18] ^ p55_add_69375_comb[13:0], p55_add_69375_comb[12:6] ^ p55_add_69375_comb[17:11] ^ p55_add_69375_comb[31:25]} + p54_add_68893;
  assign p55_add_69403_comb = (p55_add_69375_comb & p54_add_69151 ^ ~(p55_add_69375_comb | ~p54_add_69030)) + {p55_add_69397_comb, p54_add_68652[3:0]};
  assign p55_add_69426_comb = p54_add_69267 + p55_add_69425_comb;
  assign p55_xor_69465_comb = p54_add_68652[3:0] ^ p54_add_68652[14:11] ^ p54_add_68652[31:28];
  assign p55_add_69462_comb = p54_add_68837 + p55_add_69461_comb;
  assign p55_add_69444_comb = p54_add_68208 + p55_add_69443_comb;
  assign p55_add_69404_comb = p55_add_69402_comb + p55_add_69403_comb;

  // Registers for pipe stage 55:
  reg [31:0] p55_add_69030;
  reg [31:0] p55_add_69151;
  reg [31:0] p55_add_69375;
  reg [31:0] p55_add_68937;
  reg [31:0] p55_add_69056;
  reg [31:0] p55_add_69174;
  reg [31:0] p55_and_69421;
  reg [31:0] p55_concat_69272;
  reg [31:0] p55_add_69426;
  reg [3:0] p55_xor_69465;
  reg [31:0] p55_add_69324;
  reg [31:0] p55_add_68972;
  reg [31:0] p55_add_69462;
  reg [31:0] p55_add_68820;
  reg [31:0] p55_add_69307;
  reg [31:0] p55_add_68669;
  reg [31:0] p55_add_69192;
  reg [31:0] p55_add_69444;
  reg [31:0] p55_add_69074;
  reg [31:0] p55_add_69289;
  reg [31:0] p55_add_68955;
  reg [31:0] p55_add_68803;
  reg [31:0] p55_add_68438;
  reg [31:0] p55_add_69404;
  reg [31:0] p55_add_68652;
  reg [31:0] p55_add_68325;
  always_ff @ (posedge clk) begin
    p55_add_69030 <= p54_add_69030;
    p55_add_69151 <= p54_add_69151;
    p55_add_69375 <= p55_add_69375_comb;
    p55_add_68937 <= p54_add_68937;
    p55_add_69056 <= p54_add_69056;
    p55_add_69174 <= p54_add_69174;
    p55_and_69421 <= p55_and_69421_comb;
    p55_concat_69272 <= p54_concat_69272;
    p55_add_69426 <= p55_add_69426_comb;
    p55_xor_69465 <= p55_xor_69465_comb;
    p55_add_69324 <= p54_add_69324;
    p55_add_68972 <= p54_add_68972;
    p55_add_69462 <= p55_add_69462_comb;
    p55_add_68820 <= p54_add_68820;
    p55_add_69307 <= p54_add_69307;
    p55_add_68669 <= p54_add_68669;
    p55_add_69192 <= p54_add_69192;
    p55_add_69444 <= p55_add_69444_comb;
    p55_add_69074 <= p54_add_69074;
    p55_add_69289 <= p54_add_69289;
    p55_add_68955 <= p54_add_68955;
    p55_add_68803 <= p54_add_68803;
    p55_add_68438 <= p54_add_68438;
    p55_add_69404 <= p55_add_69404_comb;
    p55_add_68652 <= p54_add_68652;
    p55_add_68325 <= p54_add_68325;
  end

  // ===== Pipe stage 56:
  wire [31:0] p56_add_69518_comb;
  wire [31:0] p56_and_69569_comb;
  wire [30:0] p56_add_69540_comb;
  wire [28:0] p56_add_69550_comb;
  wire [31:0] p56_add_69573_comb;
  wire [28:0] p56_add_69595_comb;
  wire [31:0] p56_add_69614_comb;
  wire [31:0] p56_add_69591_comb;
  wire [31:0] p56_add_69545_comb;
  wire [31:0] p56_add_69546_comb;
  wire [31:0] p56_concat_69552_comb;
  wire [31:0] p56_add_69574_comb;
  wire [31:0] p56_concat_69597_comb;
  wire [31:0] p56_concat_69631_comb;
  wire [31:0] p56_add_69615_comb;
  wire [31:0] p56_add_69592_comb;
  wire [31:0] p56_add_69547_comb;
  assign p56_add_69518_comb = p55_add_68937 + p55_add_69404;
  assign p56_and_69569_comb = p55_add_69426 & p55_add_69174;
  assign p56_add_69540_comb = p55_add_68438[31:1] + 31'h0cd2_608b;
  assign p56_add_69550_comb = p55_add_68803[31:3] + 29'h03c6_ed81;
  assign p56_add_69573_comb = {p55_add_69426[1:0] ^ p55_add_69426[12:11] ^ p55_add_69426[21:20], p55_add_69426[31:21] ^ p55_add_69426[10:0] ^ p55_add_69426[19:9], p55_add_69426[20:12] ^ p55_add_69426[31:23] ^ p55_add_69426[8:0], p55_add_69426[11:2] ^ p55_add_69426[22:13] ^ p55_add_69426[31:22]} + (p56_and_69569_comb ^ p55_add_69426 & p55_add_69056 ^ p55_and_69421);
  assign p56_add_69595_comb = p55_add_69462[31:3] + 29'h1198_e041;
  assign p56_add_69614_comb = p55_add_69444 + {p55_add_69462[16:7] ^ p55_add_69462[18:9], p55_add_69462[6:0] ^ p55_add_69462[8:2] ^ p55_add_69462[31:25], p55_add_69462[31:30] ^ p55_add_69462[1:0] ^ p55_add_69462[24:23], p55_add_69462[29:17] ^ p55_add_69462[31:19] ^ p55_add_69462[22:10]};
  assign p56_add_69591_comb = p55_add_68803 + {p55_add_69444[16:7] ^ p55_add_69444[18:9], p55_add_69444[6:0] ^ p55_add_69444[8:2] ^ p55_add_69444[31:25], p55_add_69444[31:30] ^ p55_add_69444[1:0] ^ p55_add_69444[24:23], p55_add_69444[29:17] ^ p55_add_69444[31:19] ^ p55_add_69444[22:10]};
  assign p56_add_69545_comb = {p56_add_69518_comb[5:0] ^ p56_add_69518_comb[10:5] ^ p56_add_69518_comb[24:19], p56_add_69518_comb[31:27] ^ p56_add_69518_comb[4:0] ^ p56_add_69518_comb[18:14], p56_add_69518_comb[26:13] ^ p56_add_69518_comb[31:18] ^ p56_add_69518_comb[13:0], p56_add_69518_comb[12:6] ^ p56_add_69518_comb[17:11] ^ p56_add_69518_comb[31:25]} + p55_add_69030;
  assign p56_add_69546_comb = (p56_add_69518_comb & p55_add_69375 ^ ~(p56_add_69518_comb | ~p55_add_69151)) + {p56_add_69540_comb, p55_add_68438[0]};
  assign p56_concat_69552_comb = {p56_add_69550_comb, p55_add_68803[2:0]};
  assign p56_add_69574_comb = p55_add_69404 + p56_add_69573_comb;
  assign p56_concat_69597_comb = {p56_add_69595_comb, p55_add_69462[2:0]};
  assign p56_concat_69631_comb = {p55_add_68438[6:4] ^ p55_add_68438[17:15], p55_add_68438[3:0] ^ p55_add_68438[14:11] ^ p55_add_68438[31:28], p55_add_68438[31:21] ^ p55_add_68438[10:0] ^ p55_add_68438[27:17], p55_add_68438[20:7] ^ p55_add_68438[31:18] ^ p55_add_68438[16:3]};
  assign p56_add_69615_comb = p55_add_69324 + p56_add_69614_comb;
  assign p56_add_69592_comb = p55_add_68669 + p56_add_69591_comb;
  assign p56_add_69547_comb = p56_add_69545_comb + p56_add_69546_comb;

  // Registers for pipe stage 56:
  reg [31:0] p56_add_69151;
  reg [31:0] p56_add_69375;
  reg [31:0] p56_add_69518;
  reg [31:0] p56_add_69056;
  reg [31:0] p56_concat_69552;
  reg [31:0] p56_add_69174;
  reg [31:0] p56_concat_69272;
  reg [31:0] p56_add_69426;
  reg [31:0] p56_and_69569;
  reg [31:0] p56_add_69574;
  reg [31:0] p56_concat_69597;
  reg [3:0] p56_xor_69465;
  reg [31:0] p56_concat_69631;
  reg [31:0] p56_add_69615;
  reg [31:0] p56_add_68972;
  reg [31:0] p56_add_68820;
  reg [31:0] p56_add_69307;
  reg [31:0] p56_add_69592;
  reg [31:0] p56_add_69192;
  reg [31:0] p56_add_69444;
  reg [31:0] p56_add_69074;
  reg [31:0] p56_add_69289;
  reg [31:0] p56_add_68955;
  reg [31:0] p56_add_69547;
  reg [31:0] p56_add_68652;
  reg [31:0] p56_add_68325;
  always_ff @ (posedge clk) begin
    p56_add_69151 <= p55_add_69151;
    p56_add_69375 <= p55_add_69375;
    p56_add_69518 <= p56_add_69518_comb;
    p56_add_69056 <= p55_add_69056;
    p56_concat_69552 <= p56_concat_69552_comb;
    p56_add_69174 <= p55_add_69174;
    p56_concat_69272 <= p55_concat_69272;
    p56_add_69426 <= p55_add_69426;
    p56_and_69569 <= p56_and_69569_comb;
    p56_add_69574 <= p56_add_69574_comb;
    p56_concat_69597 <= p56_concat_69597_comb;
    p56_xor_69465 <= p55_xor_69465;
    p56_concat_69631 <= p56_concat_69631_comb;
    p56_add_69615 <= p56_add_69615_comb;
    p56_add_68972 <= p55_add_68972;
    p56_add_68820 <= p55_add_68820;
    p56_add_69307 <= p55_add_69307;
    p56_add_69592 <= p56_add_69592_comb;
    p56_add_69192 <= p55_add_69192;
    p56_add_69444 <= p55_add_69444;
    p56_add_69074 <= p55_add_69074;
    p56_add_69289 <= p55_add_69289;
    p56_add_68955 <= p55_add_68955;
    p56_add_69547 <= p56_add_69547_comb;
    p56_add_68652 <= p55_add_68652;
    p56_add_68325 <= p55_add_68325;
  end

  // ===== Pipe stage 57:
  wire [31:0] p57_add_69684_comb;
  wire [31:0] p57_and_69727_comb;
  wire [31:0] p57_add_69731_comb;
  wire [31:0] p57_add_69750_comb;
  wire [31:0] p57_add_69706_comb;
  wire [31:0] p57_add_69707_comb;
  wire [31:0] p57_not_69709_comb;
  wire [31:0] p57_add_69710_comb;
  wire [31:0] p57_add_69733_comb;
  wire [31:0] p57_add_69732_comb;
  wire [31:0] p57_add_69751_comb;
  wire [31:0] p57_add_69708_comb;
  assign p57_add_69684_comb = p56_add_69056 + p56_add_69547;
  assign p57_and_69727_comb = p56_add_69574 & p56_add_69426;
  assign p57_add_69731_comb = {p56_add_69574[1:0] ^ p56_add_69574[12:11] ^ p56_add_69574[21:20], p56_add_69574[31:21] ^ p56_add_69574[10:0] ^ p56_add_69574[19:9], p56_add_69574[20:12] ^ p56_add_69574[31:23] ^ p56_add_69574[8:0], p56_add_69574[11:2] ^ p56_add_69574[22:13] ^ p56_add_69574[31:22]} + (p57_and_69727_comb ^ p56_add_69574 & p56_add_69174 ^ p56_and_69569);
  assign p57_add_69750_comb = p56_add_68955 + {p56_add_69592[16:7] ^ p56_add_69592[18:9], p56_add_69592[6:0] ^ p56_add_69592[8:2] ^ p56_add_69592[31:25], p56_add_69592[31:30] ^ p56_add_69592[1:0] ^ p56_add_69592[24:23], p56_add_69592[29:17] ^ p56_add_69592[31:19] ^ p56_add_69592[22:10]};
  assign p57_add_69706_comb = {p57_add_69684_comb[5:0] ^ p57_add_69684_comb[10:5] ^ p57_add_69684_comb[24:19], p57_add_69684_comb[31:27] ^ p57_add_69684_comb[4:0] ^ p57_add_69684_comb[18:14], p57_add_69684_comb[26:13] ^ p57_add_69684_comb[31:18] ^ p57_add_69684_comb[13:0], p57_add_69684_comb[12:6] ^ p57_add_69684_comb[17:11] ^ p57_add_69684_comb[31:25]} + p56_add_69151;
  assign p57_add_69707_comb = (p57_add_69684_comb & p56_add_69518 ^ ~(p57_add_69684_comb | ~p56_add_69375)) + p56_concat_69552;
  assign p57_not_69709_comb = ~p56_add_69518;
  assign p57_add_69710_comb = p56_add_69518 + p56_add_68955;
  assign p57_add_69733_comb = p57_add_69684_comb + p56_add_69289;
  assign p57_add_69732_comb = p56_add_69547 + p57_add_69731_comb;
  assign p57_add_69751_comb = p56_add_68820 + p57_add_69750_comb;
  assign p57_add_69708_comb = p57_add_69706_comb + p57_add_69707_comb;

  // Registers for pipe stage 57:
  reg [31:0] p57_add_69375;
  reg [31:0] p57_add_69684;
  reg [31:0] p57_add_69174;
  reg [31:0] p57_not_69709;
  reg [31:0] p57_concat_69272;
  reg [31:0] p57_add_69426;
  reg [31:0] p57_add_69710;
  reg [31:0] p57_add_69574;
  reg [31:0] p57_and_69727;
  reg [31:0] p57_add_69733;
  reg [31:0] p57_add_69732;
  reg [31:0] p57_concat_69597;
  reg [3:0] p57_xor_69465;
  reg [31:0] p57_concat_69631;
  reg [31:0] p57_add_69615;
  reg [31:0] p57_add_68972;
  reg [31:0] p57_add_69751;
  reg [31:0] p57_add_69307;
  reg [31:0] p57_add_69592;
  reg [31:0] p57_add_69192;
  reg [31:0] p57_add_69444;
  reg [31:0] p57_add_69074;
  reg [31:0] p57_add_69708;
  reg [31:0] p57_add_68652;
  reg [31:0] p57_add_68325;
  always_ff @ (posedge clk) begin
    p57_add_69375 <= p56_add_69375;
    p57_add_69684 <= p57_add_69684_comb;
    p57_add_69174 <= p56_add_69174;
    p57_not_69709 <= p57_not_69709_comb;
    p57_concat_69272 <= p56_concat_69272;
    p57_add_69426 <= p56_add_69426;
    p57_add_69710 <= p57_add_69710_comb;
    p57_add_69574 <= p56_add_69574;
    p57_and_69727 <= p57_and_69727_comb;
    p57_add_69733 <= p57_add_69733_comb;
    p57_add_69732 <= p57_add_69732_comb;
    p57_concat_69597 <= p56_concat_69597;
    p57_xor_69465 <= p56_xor_69465;
    p57_concat_69631 <= p56_concat_69631;
    p57_add_69615 <= p56_add_69615;
    p57_add_68972 <= p56_add_68972;
    p57_add_69751 <= p57_add_69751_comb;
    p57_add_69307 <= p56_add_69307;
    p57_add_69592 <= p56_add_69592;
    p57_add_69192 <= p56_add_69192;
    p57_add_69444 <= p56_add_69444;
    p57_add_69074 <= p56_add_69074;
    p57_add_69708 <= p57_add_69708_comb;
    p57_add_68652 <= p56_add_68652;
    p57_add_68325 <= p56_add_68325;
  end

  // ===== Pipe stage 58:
  wire [31:0] p58_add_69802_comb;
  wire [31:0] p58_and_69843_comb;
  wire [30:0] p58_add_69850_comb;
  wire [31:0] p58_add_69849_comb;
  wire [29:0] p58_add_69856_comb;
  wire [31:0] p58_add_69874_comb;
  wire [31:0] p58_add_69823_comb;
  wire [31:0] p58_add_69824_comb;
  wire [31:0] p58_not_69826_comb;
  wire [31:0] p58_concat_69853_comb;
  wire [31:0] p58_add_69852_comb;
  wire [31:0] p58_concat_69858_comb;
  wire [31:0] p58_add_69875_comb;
  wire [31:0] p58_add_69825_comb;
  assign p58_add_69802_comb = p57_add_69174 + p57_add_69708;
  assign p58_and_69843_comb = p57_add_69732 & p57_add_69574;
  assign p58_add_69850_comb = p57_add_69074[31:1] + 31'h276c_5525;
  assign p58_add_69849_comb = {p57_add_69732[1:0] ^ p57_add_69732[12:11] ^ p57_add_69732[21:20], p57_add_69732[31:21] ^ p57_add_69732[10:0] ^ p57_add_69732[19:9], p57_add_69732[20:12] ^ p57_add_69732[31:23] ^ p57_add_69732[8:0], p57_add_69732[11:2] ^ p57_add_69732[22:13] ^ p57_add_69732[31:22]} + (p58_and_69843_comb ^ p57_add_69732 & p57_add_69426 ^ p57_and_69727);
  assign p58_add_69856_comb = p57_add_69751[31:2] + 30'h2132_1e05;
  assign p58_add_69874_comb = p57_add_69074 + {p57_add_69751[16:7] ^ p57_add_69751[18:9], p57_add_69751[6:0] ^ p57_add_69751[8:2] ^ p57_add_69751[31:25], p57_add_69751[31:30] ^ p57_add_69751[1:0] ^ p57_add_69751[24:23], p57_add_69751[29:17] ^ p57_add_69751[31:19] ^ p57_add_69751[22:10]};
  assign p58_add_69823_comb = {p58_add_69802_comb[5:0] ^ p58_add_69802_comb[10:5] ^ p58_add_69802_comb[24:19], p58_add_69802_comb[31:27] ^ p58_add_69802_comb[4:0] ^ p58_add_69802_comb[18:14], p58_add_69802_comb[26:13] ^ p58_add_69802_comb[31:18] ^ p58_add_69802_comb[13:0], p58_add_69802_comb[12:6] ^ p58_add_69802_comb[17:11] ^ p58_add_69802_comb[31:25]} + p57_add_69375;
  assign p58_add_69824_comb = (p58_add_69802_comb & p57_add_69684 ^ ~(p58_add_69802_comb | p57_not_69709)) + p57_concat_69272;
  assign p58_not_69826_comb = ~p57_add_69684;
  assign p58_concat_69853_comb = {p58_add_69850_comb, p57_add_69074[0]};
  assign p58_add_69852_comb = p57_add_69708 + p58_add_69849_comb;
  assign p58_concat_69858_comb = {p58_add_69856_comb, p57_add_69751[1:0]};
  assign p58_add_69875_comb = p57_add_68972 + p58_add_69874_comb;
  assign p58_add_69825_comb = p58_add_69823_comb + p58_add_69824_comb;

  // Registers for pipe stage 58:
  reg [31:0] p58_add_69802;
  reg [31:0] p58_add_69426;
  reg [31:0] p58_not_69826;
  reg [31:0] p58_add_69710;
  reg [31:0] p58_add_69574;
  reg [31:0] p58_add_69733;
  reg [31:0] p58_add_69732;
  reg [31:0] p58_and_69843;
  reg [31:0] p58_concat_69853;
  reg [31:0] p58_add_69852;
  reg [31:0] p58_concat_69858;
  reg [31:0] p58_concat_69597;
  reg [3:0] p58_xor_69465;
  reg [31:0] p58_concat_69631;
  reg [31:0] p58_add_69615;
  reg [31:0] p58_add_69875;
  reg [31:0] p58_add_69307;
  reg [31:0] p58_add_69592;
  reg [31:0] p58_add_69192;
  reg [31:0] p58_add_69444;
  reg [31:0] p58_add_69825;
  reg [31:0] p58_add_68652;
  reg [31:0] p58_add_68325;
  always_ff @ (posedge clk) begin
    p58_add_69802 <= p58_add_69802_comb;
    p58_add_69426 <= p57_add_69426;
    p58_not_69826 <= p58_not_69826_comb;
    p58_add_69710 <= p57_add_69710;
    p58_add_69574 <= p57_add_69574;
    p58_add_69733 <= p57_add_69733;
    p58_add_69732 <= p57_add_69732;
    p58_and_69843 <= p58_and_69843_comb;
    p58_concat_69853 <= p58_concat_69853_comb;
    p58_add_69852 <= p58_add_69852_comb;
    p58_concat_69858 <= p58_concat_69858_comb;
    p58_concat_69597 <= p57_concat_69597;
    p58_xor_69465 <= p57_xor_69465;
    p58_concat_69631 <= p57_concat_69631;
    p58_add_69615 <= p57_add_69615;
    p58_add_69875 <= p58_add_69875_comb;
    p58_add_69307 <= p57_add_69307;
    p58_add_69592 <= p57_add_69592;
    p58_add_69192 <= p57_add_69192;
    p58_add_69444 <= p57_add_69444;
    p58_add_69825 <= p58_add_69825_comb;
    p58_add_68652 <= p57_add_68652;
    p58_add_68325 <= p57_add_68325;
  end

  // ===== Pipe stage 59:
  wire [31:0] p59_add_69922_comb;
  wire [31:0] p59_and_69962_comb;
  wire [31:0] p59_add_69966_comb;
  wire [31:0] p59_add_69943_comb;
  wire [31:0] p59_add_69967_comb;
  wire [31:0] p59_add_69968_comb;
  wire [31:0] p59_add_69945_comb;
  assign p59_add_69922_comb = p58_add_69426 + p58_add_69825;
  assign p59_and_69962_comb = p58_add_69852 & p58_add_69732;
  assign p59_add_69966_comb = {p58_add_69852[1:0] ^ p58_add_69852[12:11] ^ p58_add_69852[21:20], p58_add_69852[31:21] ^ p58_add_69852[10:0] ^ p58_add_69852[19:9], p58_add_69852[20:12] ^ p58_add_69852[31:23] ^ p58_add_69852[8:0], p58_add_69852[11:2] ^ p58_add_69852[22:13] ^ p58_add_69852[31:22]} + (p59_and_69962_comb ^ p58_add_69852 & p58_add_69574 ^ p58_and_69843);
  assign p59_add_69943_comb = {p59_add_69922_comb[5:0] ^ p59_add_69922_comb[10:5] ^ p59_add_69922_comb[24:19], p59_add_69922_comb[31:27] ^ p59_add_69922_comb[4:0] ^ p59_add_69922_comb[18:14], p59_add_69922_comb[26:13] ^ p59_add_69922_comb[31:18] ^ p59_add_69922_comb[13:0], p59_add_69922_comb[12:6] ^ p59_add_69922_comb[17:11] ^ p59_add_69922_comb[31:25]} + (p59_add_69922_comb & p58_add_69802 ^ ~(p59_add_69922_comb | p58_not_69826));
  assign p59_add_69967_comb = p58_add_69825 + p59_add_69966_comb;
  assign p59_add_69968_comb = p59_add_69922_comb + p58_add_69444;
  assign p59_add_69945_comb = p59_add_69943_comb + 32'h34b0_bcb5;

  // Registers for pipe stage 59:
  reg [31:0] p59_add_69802;
  reg [31:0] p59_add_69922;
  reg [31:0] p59_add_69710;
  reg [31:0] p59_add_69574;
  reg [31:0] p59_add_69733;
  reg [31:0] p59_add_69732;
  reg [31:0] p59_concat_69853;
  reg [31:0] p59_add_69852;
  reg [31:0] p59_and_69962;
  reg [31:0] p59_add_69967;
  reg [31:0] p59_add_69968;
  reg [31:0] p59_concat_69858;
  reg [31:0] p59_concat_69597;
  reg [3:0] p59_xor_69465;
  reg [31:0] p59_concat_69631;
  reg [31:0] p59_add_69945;
  reg [31:0] p59_add_69615;
  reg [31:0] p59_add_69875;
  reg [31:0] p59_add_69307;
  reg [31:0] p59_add_69592;
  reg [31:0] p59_add_69192;
  reg [31:0] p59_add_68652;
  reg [31:0] p59_add_68325;
  always_ff @ (posedge clk) begin
    p59_add_69802 <= p58_add_69802;
    p59_add_69922 <= p59_add_69922_comb;
    p59_add_69710 <= p58_add_69710;
    p59_add_69574 <= p58_add_69574;
    p59_add_69733 <= p58_add_69733;
    p59_add_69732 <= p58_add_69732;
    p59_concat_69853 <= p58_concat_69853;
    p59_add_69852 <= p58_add_69852;
    p59_and_69962 <= p59_and_69962_comb;
    p59_add_69967 <= p59_add_69967_comb;
    p59_add_69968 <= p59_add_69968_comb;
    p59_concat_69858 <= p58_concat_69858;
    p59_concat_69597 <= p58_concat_69597;
    p59_xor_69465 <= p58_xor_69465;
    p59_concat_69631 <= p58_concat_69631;
    p59_add_69945 <= p59_add_69945_comb;
    p59_add_69615 <= p58_add_69615;
    p59_add_69875 <= p58_add_69875;
    p59_add_69307 <= p58_add_69307;
    p59_add_69592 <= p58_add_69592;
    p59_add_69192 <= p58_add_69192;
    p59_add_68652 <= p58_add_68652;
    p59_add_68325 <= p58_add_68325;
  end

  // ===== Pipe stage 60:
  wire [31:0] p60_add_70015_comb;
  wire [31:0] p60_add_70016_comb;
  wire [31:0] p60_and_70056_comb;
  wire [31:0] p60_add_70060_comb;
  wire [31:0] p60_add_70038_comb;
  wire [31:0] p60_not_70039_comb;
  wire [31:0] p60_add_70061_comb;
  assign p60_add_70015_comb = p59_add_69945 + p59_add_69710;
  assign p60_add_70016_comb = p59_add_69574 + p60_add_70015_comb;
  assign p60_and_70056_comb = p59_add_69967 & p59_add_69852;
  assign p60_add_70060_comb = {p59_add_69967[1:0] ^ p59_add_69967[12:11] ^ p59_add_69967[21:20], p59_add_69967[31:21] ^ p59_add_69967[10:0] ^ p59_add_69967[19:9], p59_add_69967[20:12] ^ p59_add_69967[31:23] ^ p59_add_69967[8:0], p59_add_69967[11:2] ^ p59_add_69967[22:13] ^ p59_add_69967[31:22]} + (p60_and_70056_comb ^ p59_add_69967 & p59_add_69732 ^ p59_and_69962);
  assign p60_add_70038_comb = {p60_add_70016_comb[5:0] ^ p60_add_70016_comb[10:5] ^ p60_add_70016_comb[24:19], p60_add_70016_comb[31:27] ^ p60_add_70016_comb[4:0] ^ p60_add_70016_comb[18:14], p60_add_70016_comb[26:13] ^ p60_add_70016_comb[31:18] ^ p60_add_70016_comb[13:0], p60_add_70016_comb[12:6] ^ p60_add_70016_comb[17:11] ^ p60_add_70016_comb[31:25]} + (p60_add_70016_comb & p59_add_69922 ^ ~(p60_add_70016_comb | ~p59_add_69802));
  assign p60_not_70039_comb = ~p59_add_69922;
  assign p60_add_70061_comb = p60_add_70015_comb + p60_add_70060_comb;

  // Registers for pipe stage 60:
  reg [31:0] p60_add_69802;
  reg [31:0] p60_add_70016;
  reg [31:0] p60_add_70038;
  reg [31:0] p60_add_69733;
  reg [31:0] p60_add_69732;
  reg [31:0] p60_not_70039;
  reg [31:0] p60_concat_69853;
  reg [31:0] p60_add_69852;
  reg [31:0] p60_add_69967;
  reg [31:0] p60_add_69968;
  reg [31:0] p60_and_70056;
  reg [31:0] p60_add_70061;
  reg [31:0] p60_concat_69858;
  reg [31:0] p60_concat_69597;
  reg [3:0] p60_xor_69465;
  reg [31:0] p60_concat_69631;
  reg [31:0] p60_add_69615;
  reg [31:0] p60_add_69875;
  reg [31:0] p60_add_69307;
  reg [31:0] p60_add_69592;
  reg [31:0] p60_add_69192;
  reg [31:0] p60_add_68652;
  reg [31:0] p60_add_68325;
  always_ff @ (posedge clk) begin
    p60_add_69802 <= p59_add_69802;
    p60_add_70016 <= p60_add_70016_comb;
    p60_add_70038 <= p60_add_70038_comb;
    p60_add_69733 <= p59_add_69733;
    p60_add_69732 <= p59_add_69732;
    p60_not_70039 <= p60_not_70039_comb;
    p60_concat_69853 <= p59_concat_69853;
    p60_add_69852 <= p59_add_69852;
    p60_add_69967 <= p59_add_69967;
    p60_add_69968 <= p59_add_69968;
    p60_and_70056 <= p60_and_70056_comb;
    p60_add_70061 <= p60_add_70061_comb;
    p60_concat_69858 <= p59_concat_69858;
    p60_concat_69597 <= p59_concat_69597;
    p60_xor_69465 <= p59_xor_69465;
    p60_concat_69631 <= p59_concat_69631;
    p60_add_69615 <= p59_add_69615;
    p60_add_69875 <= p59_add_69875;
    p60_add_69307 <= p59_add_69307;
    p60_add_69592 <= p59_add_69592;
    p60_add_69192 <= p59_add_69192;
    p60_add_68652 <= p59_add_68652;
    p60_add_68325 <= p59_add_68325;
  end

  // ===== Pipe stage 61:
  wire [31:0] p61_add_70109_comb;
  wire [31:0] p61_add_70110_comb;
  wire [31:0] p61_and_70131_comb;
  wire [31:0] p61_add_70111_comb;
  wire [31:0] p61_add_70135_comb;
  wire [31:0] p61_xor_70114_comb;
  wire [31:0] p61_add_70136_comb;
  assign p61_add_70109_comb = p60_add_70038 + 32'h391c_0cb3;
  assign p61_add_70110_comb = p61_add_70109_comb + p60_add_69733;
  assign p61_and_70131_comb = p60_add_70061 & p60_add_69967;
  assign p61_add_70111_comb = p60_add_69732 + p61_add_70110_comb;
  assign p61_add_70135_comb = {p60_add_70061[1:0] ^ p60_add_70061[12:11] ^ p60_add_70061[21:20], p60_add_70061[31:21] ^ p60_add_70061[10:0] ^ p60_add_70061[19:9], p60_add_70061[20:12] ^ p60_add_70061[31:23] ^ p60_add_70061[8:0], p60_add_70061[11:2] ^ p60_add_70061[22:13] ^ p60_add_70061[31:22]} + (p61_and_70131_comb ^ p60_add_70061 & p60_add_69852 ^ p60_and_70056);
  assign p61_xor_70114_comb = p61_add_70111_comb & p60_add_70016 ^ ~(p61_add_70111_comb | p60_not_70039);
  assign p61_add_70136_comb = p61_add_70110_comb + p61_add_70135_comb;

  // Registers for pipe stage 61:
  reg [31:0] p61_add_69802;
  reg [31:0] p61_add_70016;
  reg [31:0] p61_add_70111;
  reg [31:0] p61_xor_70114;
  reg [31:0] p61_concat_69853;
  reg [31:0] p61_add_69852;
  reg [31:0] p61_add_69967;
  reg [31:0] p61_add_69968;
  reg [31:0] p61_add_70061;
  reg [31:0] p61_and_70131;
  reg [31:0] p61_add_70136;
  reg [31:0] p61_concat_69858;
  reg [31:0] p61_concat_69597;
  reg [3:0] p61_xor_69465;
  reg [31:0] p61_concat_69631;
  reg [31:0] p61_add_69615;
  reg [31:0] p61_add_69875;
  reg [31:0] p61_add_69307;
  reg [31:0] p61_add_69592;
  reg [31:0] p61_add_69192;
  reg [31:0] p61_add_68652;
  reg [31:0] p61_add_68325;
  always_ff @ (posedge clk) begin
    p61_add_69802 <= p60_add_69802;
    p61_add_70016 <= p60_add_70016;
    p61_add_70111 <= p61_add_70111_comb;
    p61_xor_70114 <= p61_xor_70114_comb;
    p61_concat_69853 <= p60_concat_69853;
    p61_add_69852 <= p60_add_69852;
    p61_add_69967 <= p60_add_69967;
    p61_add_69968 <= p60_add_69968;
    p61_add_70061 <= p60_add_70061;
    p61_and_70131 <= p61_and_70131_comb;
    p61_add_70136 <= p61_add_70136_comb;
    p61_concat_69858 <= p60_concat_69858;
    p61_concat_69597 <= p60_concat_69597;
    p61_xor_69465 <= p60_xor_69465;
    p61_concat_69631 <= p60_concat_69631;
    p61_add_69615 <= p60_add_69615;
    p61_add_69875 <= p60_add_69875;
    p61_add_69307 <= p60_add_69307;
    p61_add_69592 <= p60_add_69592;
    p61_add_69192 <= p60_add_69192;
    p61_add_68652 <= p60_add_68652;
    p61_add_68325 <= p60_add_68325;
  end

  // ===== Pipe stage 62:
  wire [31:0] p62_and_70218_comb;
  wire [31:0] p62_add_70198_comb;
  wire [31:0] p62_add_70199_comb;
  wire [31:0] p62_add_70200_comb;
  wire [31:0] p62_add_70222_comb;
  wire [31:0] p62_add_70201_comb;
  wire [31:0] p62_add_70223_comb;
  assign p62_and_70218_comb = p61_add_70136 & p61_add_70061;
  assign p62_add_70198_comb = {p61_add_70111[5:0] ^ p61_add_70111[10:5] ^ p61_add_70111[24:19], p61_add_70111[31:27] ^ p61_add_70111[4:0] ^ p61_add_70111[18:14], p61_add_70111[26:13] ^ p61_add_70111[31:18] ^ p61_add_70111[13:0], p61_add_70111[12:6] ^ p61_add_70111[17:11] ^ p61_add_70111[31:25]} + p61_add_69802;
  assign p62_add_70199_comb = p61_xor_70114 + p61_concat_69853;
  assign p62_add_70200_comb = p62_add_70198_comb + p62_add_70199_comb;
  assign p62_add_70222_comb = {p61_add_70136[1:0] ^ p61_add_70136[12:11] ^ p61_add_70136[21:20], p61_add_70136[31:21] ^ p61_add_70136[10:0] ^ p61_add_70136[19:9], p61_add_70136[20:12] ^ p61_add_70136[31:23] ^ p61_add_70136[8:0], p61_add_70136[11:2] ^ p61_add_70136[22:13] ^ p61_add_70136[31:22]} + (p62_and_70218_comb ^ p61_add_70136 & p61_add_69967 ^ p61_and_70131);
  assign p62_add_70201_comb = p61_add_69852 + p62_add_70200_comb;
  assign p62_add_70223_comb = p62_add_70200_comb + p62_add_70222_comb;

  // Registers for pipe stage 62:
  reg [31:0] p62_add_70016;
  reg [31:0] p62_add_70111;
  reg [31:0] p62_add_70201;
  reg [31:0] p62_add_69967;
  reg [31:0] p62_add_69968;
  reg [31:0] p62_add_70061;
  reg [31:0] p62_add_70136;
  reg [31:0] p62_and_70218;
  reg [31:0] p62_add_70223;
  reg [31:0] p62_concat_69858;
  reg [31:0] p62_concat_69597;
  reg [3:0] p62_xor_69465;
  reg [31:0] p62_concat_69631;
  reg [31:0] p62_add_69615;
  reg [31:0] p62_add_69875;
  reg [31:0] p62_add_69307;
  reg [31:0] p62_add_69592;
  reg [31:0] p62_add_69192;
  reg [31:0] p62_add_68652;
  reg [31:0] p62_add_68325;
  always_ff @ (posedge clk) begin
    p62_add_70016 <= p61_add_70016;
    p62_add_70111 <= p61_add_70111;
    p62_add_70201 <= p62_add_70201_comb;
    p62_add_69967 <= p61_add_69967;
    p62_add_69968 <= p61_add_69968;
    p62_add_70061 <= p61_add_70061;
    p62_add_70136 <= p61_add_70136;
    p62_and_70218 <= p62_and_70218_comb;
    p62_add_70223 <= p62_add_70223_comb;
    p62_concat_69858 <= p61_concat_69858;
    p62_concat_69597 <= p61_concat_69597;
    p62_xor_69465 <= p61_xor_69465;
    p62_concat_69631 <= p61_concat_69631;
    p62_add_69615 <= p61_add_69615;
    p62_add_69875 <= p61_add_69875;
    p62_add_69307 <= p61_add_69307;
    p62_add_69592 <= p61_add_69592;
    p62_add_69192 <= p61_add_69192;
    p62_add_68652 <= p61_add_68652;
    p62_add_68325 <= p61_add_68325;
  end

  // ===== Pipe stage 63:
  wire [31:0] p63_add_70285_comb;
  wire [31:0] p63_add_70287_comb;
  wire [31:0] p63_add_70288_comb;
  wire [31:0] p63_add_70289_comb;
  wire [31:0] p63_add_70290_comb;
  assign p63_add_70285_comb = {p62_add_70201[5:0] ^ p62_add_70201[10:5] ^ p62_add_70201[24:19], p62_add_70201[31:27] ^ p62_add_70201[4:0] ^ p62_add_70201[18:14], p62_add_70201[26:13] ^ p62_add_70201[31:18] ^ p62_add_70201[13:0], p62_add_70201[12:6] ^ p62_add_70201[17:11] ^ p62_add_70201[31:25]} + (p62_add_70201 & p62_add_70111 ^ ~(p62_add_70201 | ~p62_add_70016));
  assign p63_add_70287_comb = p63_add_70285_comb + 32'h5b9c_ca4f;
  assign p63_add_70288_comb = p63_add_70287_comb + p62_add_69968;
  assign p63_add_70289_comb = p62_add_70016 + p62_add_69192;
  assign p63_add_70290_comb = p62_add_70201 + p62_add_69307;

  // Registers for pipe stage 63:
  reg [31:0] p63_add_70111;
  reg [31:0] p63_add_70201;
  reg [31:0] p63_add_69967;
  reg [31:0] p63_add_70288;
  reg [31:0] p63_add_70061;
  reg [31:0] p63_add_70289;
  reg [31:0] p63_add_70136;
  reg [31:0] p63_and_70218;
  reg [31:0] p63_add_70223;
  reg [31:0] p63_add_70290;
  reg [31:0] p63_concat_69858;
  reg [31:0] p63_concat_69597;
  reg [3:0] p63_xor_69465;
  reg [31:0] p63_concat_69631;
  reg [31:0] p63_add_69615;
  reg [31:0] p63_add_69875;
  reg [31:0] p63_add_69592;
  reg [31:0] p63_add_69192;
  reg [31:0] p63_add_68652;
  reg [31:0] p63_add_68325;
  always_ff @ (posedge clk) begin
    p63_add_70111 <= p62_add_70111;
    p63_add_70201 <= p62_add_70201;
    p63_add_69967 <= p62_add_69967;
    p63_add_70288 <= p63_add_70288_comb;
    p63_add_70061 <= p62_add_70061;
    p63_add_70289 <= p63_add_70289_comb;
    p63_add_70136 <= p62_add_70136;
    p63_and_70218 <= p62_and_70218;
    p63_add_70223 <= p62_add_70223;
    p63_add_70290 <= p63_add_70290_comb;
    p63_concat_69858 <= p62_concat_69858;
    p63_concat_69597 <= p62_concat_69597;
    p63_xor_69465 <= p62_xor_69465;
    p63_concat_69631 <= p62_concat_69631;
    p63_add_69615 <= p62_add_69615;
    p63_add_69875 <= p62_add_69875;
    p63_add_69592 <= p62_add_69592;
    p63_add_69192 <= p62_add_69192;
    p63_add_68652 <= p62_add_68652;
    p63_add_68325 <= p62_add_68325;
  end

  // ===== Pipe stage 64:
  wire [31:0] p64_add_70331_comb;
  wire [31:0] p64_and_70373_comb;
  wire [31:0] p64_add_70377_comb;
  wire [31:0] p64_add_70353_comb;
  wire [31:0] p64_not_70356_comb;
  wire [31:0] p64_add_70378_comb;
  wire [31:0] p64_add_70355_comb;
  assign p64_add_70331_comb = p63_add_69967 + p63_add_70288;
  assign p64_and_70373_comb = p63_add_70223 & p63_add_70136;
  assign p64_add_70377_comb = {p63_add_70223[1:0] ^ p63_add_70223[12:11] ^ p63_add_70223[21:20], p63_add_70223[31:21] ^ p63_add_70223[10:0] ^ p63_add_70223[19:9], p63_add_70223[20:12] ^ p63_add_70223[31:23] ^ p63_add_70223[8:0], p63_add_70223[11:2] ^ p63_add_70223[22:13] ^ p63_add_70223[31:22]} + (p64_and_70373_comb ^ p63_add_70223 & p63_add_70061 ^ p63_and_70218);
  assign p64_add_70353_comb = {p64_add_70331_comb[5:0] ^ p64_add_70331_comb[10:5] ^ p64_add_70331_comb[24:19], p64_add_70331_comb[31:27] ^ p64_add_70331_comb[4:0] ^ p64_add_70331_comb[18:14], p64_add_70331_comb[26:13] ^ p64_add_70331_comb[31:18] ^ p64_add_70331_comb[13:0], p64_add_70331_comb[12:6] ^ p64_add_70331_comb[17:11] ^ p64_add_70331_comb[31:25]} + (p64_add_70331_comb & p63_add_70201 ^ ~(p64_add_70331_comb | ~p63_add_70111));
  assign p64_not_70356_comb = ~p63_add_70201;
  assign p64_add_70378_comb = p63_add_70288 + p64_add_70377_comb;
  assign p64_add_70355_comb = p64_add_70353_comb + 32'h682e_6ff3;

  // Registers for pipe stage 64:
  reg [31:0] p64_add_70111;
  reg [31:0] p64_add_70331;
  reg [31:0] p64_add_70061;
  reg [31:0] p64_add_70289;
  reg [31:0] p64_not_70356;
  reg [31:0] p64_add_70136;
  reg [31:0] p64_add_70223;
  reg [31:0] p64_and_70373;
  reg [31:0] p64_add_70378;
  reg [31:0] p64_add_70290;
  reg [31:0] p64_concat_69858;
  reg [31:0] p64_concat_69597;
  reg [3:0] p64_xor_69465;
  reg [31:0] p64_concat_69631;
  reg [31:0] p64_add_70355;
  reg [31:0] p64_add_69615;
  reg [31:0] p64_add_69875;
  reg [31:0] p64_add_69592;
  reg [31:0] p64_add_69192;
  reg [31:0] p64_add_68652;
  reg [31:0] p64_add_68325;
  always_ff @ (posedge clk) begin
    p64_add_70111 <= p63_add_70111;
    p64_add_70331 <= p64_add_70331_comb;
    p64_add_70061 <= p63_add_70061;
    p64_add_70289 <= p63_add_70289;
    p64_not_70356 <= p64_not_70356_comb;
    p64_add_70136 <= p63_add_70136;
    p64_add_70223 <= p63_add_70223;
    p64_and_70373 <= p64_and_70373_comb;
    p64_add_70378 <= p64_add_70378_comb;
    p64_add_70290 <= p63_add_70290;
    p64_concat_69858 <= p63_concat_69858;
    p64_concat_69597 <= p63_concat_69597;
    p64_xor_69465 <= p63_xor_69465;
    p64_concat_69631 <= p63_concat_69631;
    p64_add_70355 <= p64_add_70355_comb;
    p64_add_69615 <= p63_add_69615;
    p64_add_69875 <= p63_add_69875;
    p64_add_69592 <= p63_add_69592;
    p64_add_69192 <= p63_add_69192;
    p64_add_68652 <= p63_add_68652;
    p64_add_68325 <= p63_add_68325;
  end

  // ===== Pipe stage 65:
  wire [31:0] p65_add_70421_comb;
  wire [31:0] p65_add_70422_comb;
  wire [31:0] p65_and_70466_comb;
  wire [30:0] p65_add_70443_comb;
  wire [31:0] p65_add_70470_comb;
  wire [31:0] p65_add_70471_comb;
  wire [31:0] p65_add_70448_comb;
  wire [31:0] p65_add_70449_comb;
  assign p65_add_70421_comb = p64_add_70355 + p64_add_70289;
  assign p65_add_70422_comb = p64_add_70061 + p65_add_70421_comb;
  assign p65_and_70466_comb = p64_add_70378 & p64_add_70223;
  assign p65_add_70443_comb = p64_add_69592[31:1] + 31'h3a47_c177;
  assign p65_add_70470_comb = {p64_add_70378[1:0] ^ p64_add_70378[12:11] ^ p64_add_70378[21:20], p64_add_70378[31:21] ^ p64_add_70378[10:0] ^ p64_add_70378[19:9], p64_add_70378[20:12] ^ p64_add_70378[31:23] ^ p64_add_70378[8:0], p64_add_70378[11:2] ^ p64_add_70378[22:13] ^ p64_add_70378[31:22]} + (p65_and_70466_comb ^ p64_add_70378 & p64_add_70136 ^ p64_and_70373);
  assign p65_add_70471_comb = p65_add_70421_comb + p65_add_70470_comb;
  assign p65_add_70448_comb = {p65_add_70422_comb[5:0] ^ p65_add_70422_comb[10:5] ^ p65_add_70422_comb[24:19], p65_add_70422_comb[31:27] ^ p65_add_70422_comb[4:0] ^ p65_add_70422_comb[18:14], p65_add_70422_comb[26:13] ^ p65_add_70422_comb[31:18] ^ p65_add_70422_comb[13:0], p65_add_70422_comb[12:6] ^ p65_add_70422_comb[17:11] ^ p65_add_70422_comb[31:25]} + p64_add_70111;
  assign p65_add_70449_comb = (p65_add_70422_comb & p64_add_70331 ^ ~(p65_add_70422_comb | p64_not_70356)) + {p65_add_70443_comb, p64_add_69592[0]};

  // Registers for pipe stage 65:
  reg [31:0] p65_add_70331;
  reg [31:0] p65_add_70422;
  reg [31:0] p65_add_70136;
  reg [31:0] p65_add_70223;
  reg [31:0] p65_add_70378;
  reg [31:0] p65_add_70290;
  reg [31:0] p65_and_70466;
  reg [31:0] p65_concat_69858;
  reg [31:0] p65_add_70471;
  reg [31:0] p65_concat_69597;
  reg [3:0] p65_xor_69465;
  reg [31:0] p65_concat_69631;
  reg [31:0] p65_add_69615;
  reg [31:0] p65_add_69875;
  reg [31:0] p65_add_70448;
  reg [31:0] p65_add_70449;
  reg [31:0] p65_add_69592;
  reg [31:0] p65_add_69192;
  reg [31:0] p65_add_68652;
  reg [31:0] p65_add_68325;
  always_ff @ (posedge clk) begin
    p65_add_70331 <= p64_add_70331;
    p65_add_70422 <= p65_add_70422_comb;
    p65_add_70136 <= p64_add_70136;
    p65_add_70223 <= p64_add_70223;
    p65_add_70378 <= p64_add_70378;
    p65_add_70290 <= p64_add_70290;
    p65_and_70466 <= p65_and_70466_comb;
    p65_concat_69858 <= p64_concat_69858;
    p65_add_70471 <= p65_add_70471_comb;
    p65_concat_69597 <= p64_concat_69597;
    p65_xor_69465 <= p64_xor_69465;
    p65_concat_69631 <= p64_concat_69631;
    p65_add_69615 <= p64_add_69615;
    p65_add_69875 <= p64_add_69875;
    p65_add_70448 <= p65_add_70448_comb;
    p65_add_70449 <= p65_add_70449_comb;
    p65_add_69592 <= p64_add_69592;
    p65_add_69192 <= p64_add_69192;
    p65_add_68652 <= p64_add_68652;
    p65_add_68325 <= p64_add_68325;
  end

  // ===== Pipe stage 66:
  wire [31:0] p66_add_70512_comb;
  wire [31:0] p66_add_70513_comb;
  wire [31:0] p66_and_70552_comb;
  wire [31:0] p66_add_70556_comb;
  wire [31:0] p66_add_70535_comb;
  wire [31:0] p66_add_70557_comb;
  assign p66_add_70512_comb = p65_add_70448 + p65_add_70449;
  assign p66_add_70513_comb = p65_add_70136 + p66_add_70512_comb;
  assign p66_and_70552_comb = p65_add_70471 & p65_add_70378;
  assign p66_add_70556_comb = {p65_add_70471[1:0] ^ p65_add_70471[12:11] ^ p65_add_70471[21:20], p65_add_70471[31:21] ^ p65_add_70471[10:0] ^ p65_add_70471[19:9], p65_add_70471[20:12] ^ p65_add_70471[31:23] ^ p65_add_70471[8:0], p65_add_70471[11:2] ^ p65_add_70471[22:13] ^ p65_add_70471[31:22]} + (p66_and_70552_comb ^ p65_add_70471 & p65_add_70223 ^ p65_and_70466);
  assign p66_add_70535_comb = {p66_add_70513_comb[5:0] ^ p66_add_70513_comb[10:5] ^ p66_add_70513_comb[24:19], p66_add_70513_comb[31:27] ^ p66_add_70513_comb[4:0] ^ p66_add_70513_comb[18:14], p66_add_70513_comb[26:13] ^ p66_add_70513_comb[31:18] ^ p66_add_70513_comb[13:0], p66_add_70513_comb[12:6] ^ p66_add_70513_comb[17:11] ^ p66_add_70513_comb[31:25]} + (p66_add_70513_comb & p65_add_70422 ^ ~(p66_add_70513_comb | ~p65_add_70331));
  assign p66_add_70557_comb = p66_add_70512_comb + p66_add_70556_comb;

  // Registers for pipe stage 66:
  reg [31:0] p66_add_70331;
  reg [31:0] p66_add_70422;
  reg [31:0] p66_add_70223;
  reg [31:0] p66_add_70513;
  reg [31:0] p66_add_70535;
  reg [31:0] p66_add_70378;
  reg [31:0] p66_add_70290;
  reg [31:0] p66_concat_69858;
  reg [31:0] p66_add_70471;
  reg [31:0] p66_and_70552;
  reg [31:0] p66_add_70557;
  reg [31:0] p66_concat_69597;
  reg [3:0] p66_xor_69465;
  reg [31:0] p66_concat_69631;
  reg [31:0] p66_add_69615;
  reg [31:0] p66_add_69875;
  reg [31:0] p66_add_69592;
  reg [31:0] p66_add_69192;
  reg [31:0] p66_add_68652;
  reg [31:0] p66_add_68325;
  always_ff @ (posedge clk) begin
    p66_add_70331 <= p65_add_70331;
    p66_add_70422 <= p65_add_70422;
    p66_add_70223 <= p65_add_70223;
    p66_add_70513 <= p66_add_70513_comb;
    p66_add_70535 <= p66_add_70535_comb;
    p66_add_70378 <= p65_add_70378;
    p66_add_70290 <= p65_add_70290;
    p66_concat_69858 <= p65_concat_69858;
    p66_add_70471 <= p65_add_70471;
    p66_and_70552 <= p66_and_70552_comb;
    p66_add_70557 <= p66_add_70557_comb;
    p66_concat_69597 <= p65_concat_69597;
    p66_xor_69465 <= p65_xor_69465;
    p66_concat_69631 <= p65_concat_69631;
    p66_add_69615 <= p65_add_69615;
    p66_add_69875 <= p65_add_69875;
    p66_add_69592 <= p65_add_69592;
    p66_add_69192 <= p65_add_69192;
    p66_add_68652 <= p65_add_68652;
    p66_add_68325 <= p65_add_68325;
  end

  // ===== Pipe stage 67:
  wire [31:0] p67_and_70618_comb;
  wire [31:0] p67_add_70599_comb;
  wire [31:0] p67_add_70600_comb;
  wire [31:0] p67_add_70622_comb;
  wire [31:0] p67_add_70601_comb;
  wire [31:0] p67_add_70623_comb;
  assign p67_and_70618_comb = p66_add_70557 & p66_add_70471;
  assign p67_add_70599_comb = p66_add_70535 + 32'h78a5_636f;
  assign p67_add_70600_comb = p67_add_70599_comb + p66_add_70290;
  assign p67_add_70622_comb = {p66_add_70557[1:0] ^ p66_add_70557[12:11] ^ p66_add_70557[21:20], p66_add_70557[31:21] ^ p66_add_70557[10:0] ^ p66_add_70557[19:9], p66_add_70557[20:12] ^ p66_add_70557[31:23] ^ p66_add_70557[8:0], p66_add_70557[11:2] ^ p66_add_70557[22:13] ^ p66_add_70557[31:22]} + (p67_and_70618_comb ^ p66_add_70557 & p66_add_70378 ^ p66_and_70552);
  assign p67_add_70601_comb = p66_add_70223 + p67_add_70600_comb;
  assign p67_add_70623_comb = p67_add_70600_comb + p67_add_70622_comb;

  // Registers for pipe stage 67:
  reg [31:0] p67_add_70331;
  reg [31:0] p67_add_70422;
  reg [31:0] p67_add_70513;
  reg [31:0] p67_add_70378;
  reg [31:0] p67_add_70601;
  reg [31:0] p67_concat_69858;
  reg [31:0] p67_add_70471;
  reg [31:0] p67_add_70557;
  reg [31:0] p67_concat_69597;
  reg [31:0] p67_and_70618;
  reg [31:0] p67_add_70623;
  reg [3:0] p67_xor_69465;
  reg [31:0] p67_concat_69631;
  reg [31:0] p67_add_69615;
  reg [31:0] p67_add_69875;
  reg [31:0] p67_add_69592;
  reg [31:0] p67_add_69192;
  reg [31:0] p67_add_68652;
  reg [31:0] p67_add_68325;
  always_ff @ (posedge clk) begin
    p67_add_70331 <= p66_add_70331;
    p67_add_70422 <= p66_add_70422;
    p67_add_70513 <= p66_add_70513;
    p67_add_70378 <= p66_add_70378;
    p67_add_70601 <= p67_add_70601_comb;
    p67_concat_69858 <= p66_concat_69858;
    p67_add_70471 <= p66_add_70471;
    p67_add_70557 <= p66_add_70557;
    p67_concat_69597 <= p66_concat_69597;
    p67_and_70618 <= p67_and_70618_comb;
    p67_add_70623 <= p67_add_70623_comb;
    p67_xor_69465 <= p66_xor_69465;
    p67_concat_69631 <= p66_concat_69631;
    p67_add_69615 <= p66_add_69615;
    p67_add_69875 <= p66_add_69875;
    p67_add_69592 <= p66_add_69592;
    p67_add_69192 <= p66_add_69192;
    p67_add_68652 <= p66_add_68652;
    p67_add_68325 <= p66_add_68325;
  end

  // ===== Pipe stage 68:
  wire [31:0] p68_and_70703_comb;
  wire [31:0] p68_add_70683_comb;
  wire [31:0] p68_add_70684_comb;
  wire [31:0] p68_add_70685_comb;
  wire [31:0] p68_add_70707_comb;
  wire [31:0] p68_add_70686_comb;
  wire [31:0] p68_add_70708_comb;
  assign p68_and_70703_comb = p67_add_70623 & p67_add_70557;
  assign p68_add_70683_comb = {p67_add_70601[5:0] ^ p67_add_70601[10:5] ^ p67_add_70601[24:19], p67_add_70601[31:27] ^ p67_add_70601[4:0] ^ p67_add_70601[18:14], p67_add_70601[26:13] ^ p67_add_70601[31:18] ^ p67_add_70601[13:0], p67_add_70601[12:6] ^ p67_add_70601[17:11] ^ p67_add_70601[31:25]} + p67_add_70331;
  assign p68_add_70684_comb = (p67_add_70601 & p67_add_70513 ^ ~(p67_add_70601 | ~p67_add_70422)) + p67_concat_69858;
  assign p68_add_70685_comb = p68_add_70683_comb + p68_add_70684_comb;
  assign p68_add_70707_comb = {p67_add_70623[1:0] ^ p67_add_70623[12:11] ^ p67_add_70623[21:20], p67_add_70623[31:21] ^ p67_add_70623[10:0] ^ p67_add_70623[19:9], p67_add_70623[20:12] ^ p67_add_70623[31:23] ^ p67_add_70623[8:0], p67_add_70623[11:2] ^ p67_add_70623[22:13] ^ p67_add_70623[31:22]} + (p68_and_70703_comb ^ p67_add_70623 & p67_add_70471 ^ p67_and_70618);
  assign p68_add_70686_comb = p67_add_70378 + p68_add_70685_comb;
  assign p68_add_70708_comb = p68_add_70685_comb + p68_add_70707_comb;

  // Registers for pipe stage 68:
  reg [31:0] p68_add_70422;
  reg [31:0] p68_add_70513;
  reg [31:0] p68_add_70601;
  reg [31:0] p68_add_70471;
  reg [31:0] p68_add_70686;
  reg [31:0] p68_add_70557;
  reg [31:0] p68_concat_69597;
  reg [31:0] p68_add_70623;
  reg [31:0] p68_and_70703;
  reg [31:0] p68_add_70708;
  reg [3:0] p68_xor_69465;
  reg [31:0] p68_concat_69631;
  reg [31:0] p68_add_69615;
  reg [31:0] p68_add_69875;
  reg [31:0] p68_add_69592;
  reg [31:0] p68_add_69192;
  reg [31:0] p68_add_68652;
  reg [31:0] p68_add_68325;
  always_ff @ (posedge clk) begin
    p68_add_70422 <= p67_add_70422;
    p68_add_70513 <= p67_add_70513;
    p68_add_70601 <= p67_add_70601;
    p68_add_70471 <= p67_add_70471;
    p68_add_70686 <= p68_add_70686_comb;
    p68_add_70557 <= p67_add_70557;
    p68_concat_69597 <= p67_concat_69597;
    p68_add_70623 <= p67_add_70623;
    p68_and_70703 <= p68_and_70703_comb;
    p68_add_70708 <= p68_add_70708_comb;
    p68_xor_69465 <= p67_xor_69465;
    p68_concat_69631 <= p67_concat_69631;
    p68_add_69615 <= p67_add_69615;
    p68_add_69875 <= p67_add_69875;
    p68_add_69592 <= p67_add_69592;
    p68_add_69192 <= p67_add_69192;
    p68_add_68652 <= p67_add_68652;
    p68_add_68325 <= p67_add_68325;
  end

  // ===== Pipe stage 69:
  wire [31:0] p69_and_70789_comb;
  wire [31:0] p69_add_70766_comb;
  wire [31:0] p69_add_70767_comb;
  wire [31:0] p69_add_70768_comb;
  wire [31:0] p69_add_70793_comb;
  wire [31:0] p69_add_70769_comb;
  wire [30:0] p69_add_70772_comb;
  wire [31:0] p69_add_70794_comb;
  wire [31:0] p69_add_70795_comb;
  assign p69_and_70789_comb = p68_add_70708 & p68_add_70623;
  assign p69_add_70766_comb = {p68_add_70686[5:0] ^ p68_add_70686[10:5] ^ p68_add_70686[24:19], p68_add_70686[31:27] ^ p68_add_70686[4:0] ^ p68_add_70686[18:14], p68_add_70686[26:13] ^ p68_add_70686[31:18] ^ p68_add_70686[13:0], p68_add_70686[12:6] ^ p68_add_70686[17:11] ^ p68_add_70686[31:25]} + p68_add_70422;
  assign p69_add_70767_comb = (p68_add_70686 & p68_add_70601 ^ ~(p68_add_70686 | ~p68_add_70513)) + p68_concat_69597;
  assign p69_add_70768_comb = p69_add_70766_comb + p69_add_70767_comb;
  assign p69_add_70793_comb = {p68_add_70708[1:0] ^ p68_add_70708[12:11] ^ p68_add_70708[21:20], p68_add_70708[31:21] ^ p68_add_70708[10:0] ^ p68_add_70708[19:9], p68_add_70708[20:12] ^ p68_add_70708[31:23] ^ p68_add_70708[8:0], p68_add_70708[11:2] ^ p68_add_70708[22:13] ^ p68_add_70708[31:22]} + (p69_and_70789_comb ^ p68_add_70708 & p68_add_70557 ^ p68_and_70703);
  assign p69_add_70769_comb = p68_add_70471 + p69_add_70768_comb;
  assign p69_add_70772_comb = p68_add_69875[31:1] + 31'h485f_7ffd;
  assign p69_add_70794_comb = p69_add_70768_comb + p69_add_70793_comb;
  assign p69_add_70795_comb = p68_add_70686 + p68_add_69192;

  // Registers for pipe stage 69:
  reg [31:0] p69_add_70513;
  reg [31:0] p69_add_70601;
  reg [31:0] p69_add_70686;
  reg [31:0] p69_add_70557;
  reg [31:0] p69_add_70769;
  reg [31:0] p69_add_70623;
  reg [30:0] p69_add_70772;
  reg [31:0] p69_add_70708;
  reg [31:0] p69_and_70789;
  reg [31:0] p69_add_70794;
  reg [3:0] p69_xor_69465;
  reg [31:0] p69_concat_69631;
  reg [31:0] p69_add_70795;
  reg [31:0] p69_add_69615;
  reg [31:0] p69_add_69875;
  reg [31:0] p69_add_69592;
  reg [31:0] p69_add_68652;
  reg [31:0] p69_add_68325;
  always_ff @ (posedge clk) begin
    p69_add_70513 <= p68_add_70513;
    p69_add_70601 <= p68_add_70601;
    p69_add_70686 <= p68_add_70686;
    p69_add_70557 <= p68_add_70557;
    p69_add_70769 <= p69_add_70769_comb;
    p69_add_70623 <= p68_add_70623;
    p69_add_70772 <= p69_add_70772_comb;
    p69_add_70708 <= p68_add_70708;
    p69_and_70789 <= p69_and_70789_comb;
    p69_add_70794 <= p69_add_70794_comb;
    p69_xor_69465 <= p68_xor_69465;
    p69_concat_69631 <= p68_concat_69631;
    p69_add_70795 <= p69_add_70795_comb;
    p69_add_69615 <= p68_add_69615;
    p69_add_69875 <= p68_add_69875;
    p69_add_69592 <= p68_add_69592;
    p69_add_68652 <= p68_add_68652;
    p69_add_68325 <= p68_add_68325;
  end

  // ===== Pipe stage 70:
  wire [12:0] p70_xor_70913_comb;
  wire [31:0] p70_add_70855_comb;
  wire [31:0] p70_add_70856_comb;
  wire [31:0] p70_and_70877_comb;
  wire [31:0] p70_add_70857_comb;
  wire [31:0] p70_add_70858_comb;
  wire [31:0] p70_add_70882_comb;
  wire [30:0] p70_add_70920_comb;
  wire [31:0] p70_nor_70860_comb;
  wire [31:0] p70_add_70881_comb;
  wire [31:0] p70_add_70883_comb;
  wire [31:0] p70_concat_70922_comb;
  wire [31:0] p70_add_70923_comb;
  wire [31:0] p70_add_70901_comb;
  assign p70_xor_70913_comb = p69_add_69615[29:17] ^ p69_add_69615[31:19] ^ p69_add_69615[22:10];
  assign p70_add_70855_comb = {p69_add_70769[5:0] ^ p69_add_70769[10:5] ^ p69_add_70769[24:19], p69_add_70769[31:27] ^ p69_add_70769[4:0] ^ p69_add_70769[18:14], p69_add_70769[26:13] ^ p69_add_70769[31:18] ^ p69_add_70769[13:0], p69_add_70769[12:6] ^ p69_add_70769[17:11] ^ p69_add_70769[31:25]} + p69_add_70513;
  assign p70_add_70856_comb = (p69_add_70769 & p69_add_70686 ^ ~(p69_add_70769 | ~p69_add_70601)) + {p69_add_70772, p69_add_69875[0]};
  assign p70_and_70877_comb = p69_add_70794 & p69_add_70708;
  assign p70_add_70857_comb = p70_add_70855_comb + p70_add_70856_comb;
  assign p70_add_70858_comb = p69_add_70557 + p70_add_70857_comb;
  assign p70_add_70882_comb = {p69_add_70794[1:0] ^ p69_add_70794[12:11] ^ p69_add_70794[21:20], p69_add_70794[31:21] ^ p69_add_70794[10:0] ^ p69_add_70794[19:9], p69_add_70794[20:12] ^ p69_add_70794[31:23] ^ p69_add_70794[8:0], p69_add_70794[11:2] ^ p69_add_70794[22:13] ^ p69_add_70794[31:22]} + (p70_and_70877_comb ^ p69_add_70794 & p69_add_70623 ^ p69_and_70789);
  assign p70_add_70920_comb = {p69_add_69615[16:7] ^ p69_add_69615[18:9], p69_add_69615[6:0] ^ p69_add_69615[8:2] ^ p69_add_69615[31:25], p69_add_69615[31:30] ^ p69_add_69615[1:0] ^ p69_add_69615[24:23], p70_xor_70913_comb[12:1]} + 31'h6338_bc79;
  assign p70_nor_70860_comb = ~(p70_add_70858_comb | ~p69_add_70686);
  assign p70_add_70881_comb = p69_add_70601 + p69_add_69615;
  assign p70_add_70883_comb = p70_add_70857_comb + p70_add_70882_comb;
  assign p70_concat_70922_comb = {p70_add_70920_comb, p70_xor_70913_comb[0]};
  assign p70_add_70923_comb = p69_concat_69631 + p69_add_70769;
  assign p70_add_70901_comb = {p69_add_69875[16:7] ^ p69_add_69875[18:9], p69_add_69875[6:0] ^ p69_add_69875[8:2] ^ p69_add_69875[31:25], p69_add_69875[31:30] ^ p69_add_69875[1:0] ^ p69_add_69875[24:23], p69_add_69875[29:17] ^ p69_add_69875[31:19] ^ p69_add_69875[22:10]} + 32'hbef9_a3f7;

  // Registers for pipe stage 70:
  reg [31:0] p70_add_70769;
  reg [31:0] p70_add_70623;
  reg [31:0] p70_add_70708;
  reg [31:0] p70_add_70858;
  reg [31:0] p70_nor_70860;
  reg [31:0] p70_add_70794;
  reg [31:0] p70_add_70881;
  reg [31:0] p70_and_70877;
  reg [3:0] p70_xor_69465;
  reg [31:0] p70_add_70883;
  reg [31:0] p70_concat_70922;
  reg [31:0] p70_add_70923;
  reg [31:0] p70_add_70795;
  reg [31:0] p70_add_70901;
  reg [31:0] p70_add_69592;
  reg [31:0] p70_add_68652;
  reg [31:0] p70_add_68325;
  always_ff @ (posedge clk) begin
    p70_add_70769 <= p69_add_70769;
    p70_add_70623 <= p69_add_70623;
    p70_add_70708 <= p69_add_70708;
    p70_add_70858 <= p70_add_70858_comb;
    p70_nor_70860 <= p70_nor_70860_comb;
    p70_add_70794 <= p69_add_70794;
    p70_add_70881 <= p70_add_70881_comb;
    p70_and_70877 <= p70_and_70877_comb;
    p70_xor_69465 <= p69_xor_69465;
    p70_add_70883 <= p70_add_70883_comb;
    p70_concat_70922 <= p70_concat_70922_comb;
    p70_add_70923 <= p70_add_70923_comb;
    p70_add_70795 <= p69_add_70795;
    p70_add_70901 <= p70_add_70901_comb;
    p70_add_69592 <= p69_add_69592;
    p70_add_68652 <= p69_add_68652;
    p70_add_68325 <= p69_add_68325;
  end

  // ===== Pipe stage 71:
  wire [31:0] p71_add_70977_comb;
  wire [31:0] p71_add_70979_comb;
  wire [31:0] p71_add_70980_comb;
  wire [31:0] p71_not_70981_comb;
  assign p71_add_70977_comb = {p70_add_70858[5:0] ^ p70_add_70858[10:5] ^ p70_add_70858[24:19], p70_add_70858[31:27] ^ p70_add_70858[4:0] ^ p70_add_70858[18:14], p70_add_70858[26:13] ^ p70_add_70858[31:18] ^ p70_add_70858[13:0], p70_add_70858[12:6] ^ p70_add_70858[17:11] ^ p70_add_70858[31:25]} + (p70_add_70858 & p70_add_70769 ^ p70_nor_70860);
  assign p71_add_70979_comb = p71_add_70977_comb + 32'ha450_6ceb;
  assign p71_add_70980_comb = p71_add_70979_comb + p70_add_70881;
  assign p71_not_70981_comb = ~p70_add_70769;

  // Registers for pipe stage 71:
  reg [31:0] p71_add_70623;
  reg [31:0] p71_add_70708;
  reg [31:0] p71_add_70858;
  reg [31:0] p71_add_70794;
  reg [31:0] p71_add_70980;
  reg [31:0] p71_and_70877;
  reg [31:0] p71_not_70981;
  reg [3:0] p71_xor_69465;
  reg [31:0] p71_add_70883;
  reg [31:0] p71_concat_70922;
  reg [31:0] p71_add_70923;
  reg [31:0] p71_add_70795;
  reg [31:0] p71_add_70901;
  reg [31:0] p71_add_69592;
  reg [31:0] p71_add_68652;
  reg [31:0] p71_add_68325;
  always_ff @ (posedge clk) begin
    p71_add_70623 <= p70_add_70623;
    p71_add_70708 <= p70_add_70708;
    p71_add_70858 <= p70_add_70858;
    p71_add_70794 <= p70_add_70794;
    p71_add_70980 <= p71_add_70980_comb;
    p71_and_70877 <= p70_and_70877;
    p71_not_70981 <= p71_not_70981_comb;
    p71_xor_69465 <= p70_xor_69465;
    p71_add_70883 <= p70_add_70883;
    p71_concat_70922 <= p70_concat_70922;
    p71_add_70923 <= p70_add_70923;
    p71_add_70795 <= p70_add_70795;
    p71_add_70901 <= p70_add_70901;
    p71_add_69592 <= p70_add_69592;
    p71_add_68652 <= p70_add_68652;
    p71_add_68325 <= p70_add_68325;
  end

  // ===== Pipe stage 72:
  wire [31:0] p72_add_71014_comb;
  wire [31:0] p72_and_71051_comb;
  wire [31:0] p72_add_71067_comb;
  wire [31:0] p72_add_71068_comb;
  wire [31:0] p72_add_71069_comb;
  wire [31:0] p72_add_71070_comb;
  wire [31:0] p72_add_71071_comb;
  wire [31:0] p72_add_71072_comb;
  assign p72_add_71014_comb = p71_add_70623 + p71_add_70980;
  assign p72_and_71051_comb = p71_add_70883 & p71_add_70794;
  assign p72_add_71067_comb = {p71_add_70883[1:0] ^ p71_add_70883[12:11] ^ p71_add_70883[21:20], p71_add_70883[31:21] ^ p71_add_70883[10:0] ^ p71_add_70883[19:9], p71_add_70883[20:12] ^ p71_add_70883[31:23] ^ p71_add_70883[8:0], p71_add_70883[11:2] ^ p71_add_70883[22:13] ^ p71_add_70883[31:22]} + (p72_and_71051_comb ^ p71_add_70883 & p71_add_70708 ^ p71_and_70877);
  assign p72_add_71068_comb = {p72_add_71014_comb[5:0] ^ p72_add_71014_comb[10:5] ^ p72_add_71014_comb[24:19], p72_add_71014_comb[31:27] ^ p72_add_71014_comb[4:0] ^ p72_add_71014_comb[18:14], p72_add_71014_comb[26:13] ^ p72_add_71014_comb[31:18] ^ p72_add_71014_comb[13:0], p72_add_71014_comb[12:6] ^ p72_add_71014_comb[17:11] ^ p72_add_71014_comb[31:25]} + {p71_add_68652[6:4] ^ p71_add_68652[17:15], p71_xor_69465, p71_add_68652[31:21] ^ p71_add_68652[10:0] ^ p71_add_68652[27:17], p71_add_68652[20:7] ^ p71_add_68652[31:18] ^ p71_add_68652[16:3]};
  assign p72_add_71069_comb = (p72_add_71014_comb & p71_add_70858 ^ ~(p72_add_71014_comb | p71_not_70981)) + p71_add_68325;
  assign p72_add_71070_comb = p71_add_70980 + p72_add_71067_comb;
  assign p72_add_71071_comb = p71_add_70795 + p72_add_71068_comb;
  assign p72_add_71072_comb = p72_add_71069_comb + p71_add_70901;

  // Registers for pipe stage 72:
  reg [31:0] p72_add_70708;
  reg [31:0] p72_add_70858;
  reg [31:0] p72_add_70794;
  reg [31:0] p72_add_71014;
  reg [31:0] p72_add_70883;
  reg [31:0] p72_and_71051;
  reg [31:0] p72_add_71070;
  reg [31:0] p72_concat_70922;
  reg [31:0] p72_add_70923;
  reg [31:0] p72_add_71071;
  reg [31:0] p72_add_71072;
  reg [31:0] p72_add_69592;
  reg [31:0] p72_add_68652;
  always_ff @ (posedge clk) begin
    p72_add_70708 <= p71_add_70708;
    p72_add_70858 <= p71_add_70858;
    p72_add_70794 <= p71_add_70794;
    p72_add_71014 <= p72_add_71014_comb;
    p72_add_70883 <= p71_add_70883;
    p72_and_71051 <= p72_and_71051_comb;
    p72_add_71070 <= p72_add_71070_comb;
    p72_concat_70922 <= p71_concat_70922;
    p72_add_70923 <= p71_add_70923;
    p72_add_71071 <= p72_add_71071_comb;
    p72_add_71072 <= p72_add_71072_comb;
    p72_add_69592 <= p71_add_69592;
    p72_add_68652 <= p71_add_68652;
  end

  // ===== Pipe stage 73:
  wire [31:0] p73_and_71116_comb;
  wire [31:0] p73_add_71111_comb;
  wire [31:0] p73_add_71118_comb;
  wire [31:0] p73_add_71134_comb;
  wire [31:0] p73_add_71141_comb;
  wire [30:0] p73_add_71156_comb;
  wire [30:0] p73_add_71158_comb;
  wire [29:0] p73_add_71161_comb;
  wire [31:0] p73_xor_71148_comb;
  wire [31:0] p73_add_71160_comb;
  wire [31:0] p73_concat_71165_comb;
  wire [31:0] p73_concat_71166_comb;
  wire [31:0] p73_concat_71167_comb;
  wire [31:0] p73_add_71168_comb;
  wire [31:0] p73_add_71169_comb;
  wire [31:0] p73_add_71144_comb;
  wire [31:0] p73_add_71145_comb;
  assign p73_and_71116_comb = p72_add_71070 & p72_add_70883;
  assign p73_add_71111_comb = p72_add_71071 + p72_add_71072;
  assign p73_add_71118_comb = p72_add_70708 + p73_add_71111_comb;
  assign p73_add_71134_comb = {p72_add_71070[1:0] ^ p72_add_71070[12:11] ^ p72_add_71070[21:20], p72_add_71070[31:21] ^ p72_add_71070[10:0] ^ p72_add_71070[19:9], p72_add_71070[20:12] ^ p72_add_71070[31:23] ^ p72_add_71070[8:0], p72_add_71070[11:2] ^ p72_add_71070[22:13] ^ p72_add_71070[31:22]} + (p73_and_71116_comb ^ p72_add_71070 & p72_add_70794 ^ p72_and_71051);
  assign p73_add_71141_comb = p73_add_71111_comb + p73_add_71134_comb;
  assign p73_add_71156_comb = p72_add_71070[31:1] + 31'h1e37_79b9;
  assign p73_add_71158_comb = p72_add_70883[31:1] + 31'h52a7_fa9d;
  assign p73_add_71161_comb = p73_add_71118_comb[31:2] + 30'h26c1_5a23;
  assign p73_xor_71148_comb = p73_add_71141_comb & p72_add_71070 ^ p73_add_71141_comb & p72_add_70883 ^ p73_and_71116_comb;
  assign p73_add_71160_comb = p72_add_70794 + 32'h510e_527f;
  assign p73_concat_71165_comb = {p73_add_71156_comb, p72_add_71070[0]};
  assign p73_concat_71166_comb = {p73_add_71158_comb, p72_add_70883[0]};
  assign p73_concat_71167_comb = {p73_add_71161_comb, p73_add_71118_comb[1:0]};
  assign p73_add_71168_comb = p72_add_71014 + 32'h1f83_d9ab;
  assign p73_add_71169_comb = p72_add_70858 + 32'h5be0_cd19;
  assign p73_add_71144_comb = {p73_add_71118_comb[5:0] ^ p73_add_71118_comb[10:5] ^ p73_add_71118_comb[24:19], p73_add_71118_comb[31:27] ^ p73_add_71118_comb[4:0] ^ p73_add_71118_comb[18:14], p73_add_71118_comb[26:13] ^ p73_add_71118_comb[31:18] ^ p73_add_71118_comb[13:0], p73_add_71118_comb[12:6] ^ p73_add_71118_comb[17:11] ^ p73_add_71118_comb[31:25]} + p72_add_68652;
  assign p73_add_71145_comb = p72_concat_70922 + (p73_add_71118_comb & p72_add_71014 ^ ~(p73_add_71118_comb | ~p72_add_70858));

  // Registers for pipe stage 73:
  reg [31:0] p73_add_71141;
  reg [31:0] p73_xor_71148;
  reg [31:0] p73_add_71160;
  reg [31:0] p73_concat_71165;
  reg [31:0] p73_concat_71166;
  reg [31:0] p73_concat_71167;
  reg [31:0] p73_add_71168;
  reg [31:0] p73_add_71169;
  reg [31:0] p73_add_71144;
  reg [31:0] p73_add_70923;
  reg [31:0] p73_add_71145;
  reg [31:0] p73_add_69592;
  always_ff @ (posedge clk) begin
    p73_add_71141 <= p73_add_71141_comb;
    p73_xor_71148 <= p73_xor_71148_comb;
    p73_add_71160 <= p73_add_71160_comb;
    p73_concat_71165 <= p73_concat_71165_comb;
    p73_concat_71166 <= p73_concat_71166_comb;
    p73_concat_71167 <= p73_concat_71167_comb;
    p73_add_71168 <= p73_add_71168_comb;
    p73_add_71169 <= p73_add_71169_comb;
    p73_add_71144 <= p73_add_71144_comb;
    p73_add_70923 <= p72_add_70923;
    p73_add_71145 <= p73_add_71145_comb;
    p73_add_69592 <= p72_add_69592;
  end

  // ===== Pipe stage 74:
  wire [31:0] p74_add_71210_comb;
  wire [31:0] p74_add_71211_comb;
  wire [31:0] p74_add_71213_comb;
  wire [31:0] p74_add_71218_comb;
  wire [31:0] p74_add_71219_comb;
  wire [31:0] p74_add_71215_comb;
  wire [31:0] p74_add_71216_comb;
  assign p74_add_71210_comb = p73_add_71144 + p73_add_70923;
  assign p74_add_71211_comb = p73_add_71145 + p73_add_69592;
  assign p74_add_71213_comb = p74_add_71210_comb + p74_add_71211_comb;
  assign p74_add_71218_comb = p73_add_71141 + 32'hbb67_ae85;
  assign p74_add_71219_comb = p74_add_71213_comb + p73_add_71160;
  assign p74_add_71215_comb = {p73_add_71141[1:0] ^ p73_add_71141[12:11] ^ p73_add_71141[21:20], p73_add_71141[31:21] ^ p73_add_71141[10:0] ^ p73_add_71141[19:9], p73_add_71141[20:12] ^ p73_add_71141[31:23] ^ p73_add_71141[8:0], p73_add_71141[11:2] ^ p73_add_71141[22:13] ^ p73_add_71141[31:22]} + p74_add_71213_comb;
  assign p74_add_71216_comb = p73_xor_71148 + 32'h6a09_e667;

  // Registers for pipe stage 74:
  reg [31:0] p74_add_71218;
  reg [31:0] p74_concat_71165;
  reg [31:0] p74_concat_71166;
  reg [31:0] p74_add_71219;
  reg [31:0] p74_concat_71167;
  reg [31:0] p74_add_71168;
  reg [31:0] p74_add_71169;
  reg [31:0] p74_add_71215;
  reg [31:0] p74_add_71216;
  always_ff @ (posedge clk) begin
    p74_add_71218 <= p74_add_71218_comb;
    p74_concat_71165 <= p73_concat_71165;
    p74_concat_71166 <= p73_concat_71166;
    p74_add_71219 <= p74_add_71219_comb;
    p74_concat_71167 <= p73_concat_71167;
    p74_add_71168 <= p73_add_71168;
    p74_add_71169 <= p73_add_71169;
    p74_add_71215 <= p74_add_71215_comb;
    p74_add_71216 <= p74_add_71216_comb;
  end

  // ===== Pipe stage 75:
  wire [31:0] p75_add_71238_comb;
  wire [255:0] p75_tuple_71239_comb;
  assign p75_add_71238_comb = p74_add_71215 + p74_add_71216;
  assign p75_tuple_71239_comb = {p75_add_71238_comb, p74_add_71218, p74_concat_71165, p74_concat_71166, p74_add_71219, p74_concat_71167, p74_add_71168, p74_add_71169};

  // Registers for pipe stage 75:
  reg [255:0] p75_tuple_71239;
  always_ff @ (posedge clk) begin
    p75_tuple_71239 <= p75_tuple_71239_comb;
  end
  assign out = p75_tuple_71239;
endmodule
