module xls_test(
  input wire clk,
  input wire [31:0] pc,
  input wire [31:0] ins,
  input wire [1023:0] regs,
  input wire [127:0] dmem,
  output wire [1183:0] out
);
  wire [31:0] regs_unflattened[32];
  assign regs_unflattened[0] = regs[31:0];
  assign regs_unflattened[1] = regs[63:32];
  assign regs_unflattened[2] = regs[95:64];
  assign regs_unflattened[3] = regs[127:96];
  assign regs_unflattened[4] = regs[159:128];
  assign regs_unflattened[5] = regs[191:160];
  assign regs_unflattened[6] = regs[223:192];
  assign regs_unflattened[7] = regs[255:224];
  assign regs_unflattened[8] = regs[287:256];
  assign regs_unflattened[9] = regs[319:288];
  assign regs_unflattened[10] = regs[351:320];
  assign regs_unflattened[11] = regs[383:352];
  assign regs_unflattened[12] = regs[415:384];
  assign regs_unflattened[13] = regs[447:416];
  assign regs_unflattened[14] = regs[479:448];
  assign regs_unflattened[15] = regs[511:480];
  assign regs_unflattened[16] = regs[543:512];
  assign regs_unflattened[17] = regs[575:544];
  assign regs_unflattened[18] = regs[607:576];
  assign regs_unflattened[19] = regs[639:608];
  assign regs_unflattened[20] = regs[671:640];
  assign regs_unflattened[21] = regs[703:672];
  assign regs_unflattened[22] = regs[735:704];
  assign regs_unflattened[23] = regs[767:736];
  assign regs_unflattened[24] = regs[799:768];
  assign regs_unflattened[25] = regs[831:800];
  assign regs_unflattened[26] = regs[863:832];
  assign regs_unflattened[27] = regs[895:864];
  assign regs_unflattened[28] = regs[927:896];
  assign regs_unflattened[29] = regs[959:928];
  assign regs_unflattened[30] = regs[991:960];
  assign regs_unflattened[31] = regs[1023:992];
  wire [7:0] dmem_unflattened[16];
  assign dmem_unflattened[0] = dmem[7:0];
  assign dmem_unflattened[1] = dmem[15:8];
  assign dmem_unflattened[2] = dmem[23:16];
  assign dmem_unflattened[3] = dmem[31:24];
  assign dmem_unflattened[4] = dmem[39:32];
  assign dmem_unflattened[5] = dmem[47:40];
  assign dmem_unflattened[6] = dmem[55:48];
  assign dmem_unflattened[7] = dmem[63:56];
  assign dmem_unflattened[8] = dmem[71:64];
  assign dmem_unflattened[9] = dmem[79:72];
  assign dmem_unflattened[10] = dmem[87:80];
  assign dmem_unflattened[11] = dmem[95:88];
  assign dmem_unflattened[12] = dmem[103:96];
  assign dmem_unflattened[13] = dmem[111:104];
  assign dmem_unflattened[14] = dmem[119:112];
  assign dmem_unflattened[15] = dmem[127:120];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_pc;
  reg [31:0] p0_ins;
  reg [31:0] p0_regs[32];
  reg [7:0] p0_dmem[16];
  always_ff @ (posedge clk) begin
    p0_pc <= pc;
    p0_ins <= ins;
    p0_regs <= regs_unflattened;
    p0_dmem <= dmem_unflattened;
  end

  // ===== Pipe stage 1:
  wire [11:0] p1_bit_slice_3549_comb;
  wire p1_eq_3551_comb;
  wire p1_eq_3552_comb;
  wire p1_eq_3553_comb;
  wire p1_eq_3554_comb;
  wire p1_eq_3555_comb;
  wire p1_eq_3556_comb;
  wire [31:0] p1_concat_3557_comb;
  wire [31:0] p1_array_index_3558_comb;
  wire [6:0] p1_concat_3561_comb;
  wire [31:0] p1_add_3564_comb;
  wire p1_eq_3569_comb;
  wire p1_eq_3577_comb;
  wire p1_eq_3571_comb;
  wire [7:0] p1_one_hot_3570_comb;
  wire p1_eq_3572_comb;
  wire p1_eq_3594_comb;
  wire p1_eq_3595_comb;
  wire p1_or_3596_comb;
  wire p1_eq_3597_comb;
  wire p1_eq_3598_comb;
  wire p1_eq_3599_comb;
  wire [30:0] p1_add_3587_comb;
  wire [11:0] p1_concat_3612_comb;
  wire p1_or_3615_comb;
  wire [12:0] p1_concat_3629_comb;
  wire [31:0] p1_array_index_3631_comb;
  wire [1:0] p1_concat_3601_comb;
  wire [6:0] p1_and_3602_comb;
  wire [4:0] p1_and_3604_comb;
  wire p1_and_3637_comb;
  wire p1_ugt_3667_comb;
  wire [31:0] p1_concat_3668_comb;
  wire [12:0] p1_add_3670_comb;
  wire [1:0] p1_and_3616_comb;
  wire [7:0] p1_array_index_3619_comb;
  wire [31:0] p1_add_3620_comb;
  wire [7:0] p1_array_index_3623_comb;
  wire [31:0] p1_add_3624_comb;
  wire [29:0] p1_add_3626_comb;
  wire [30:0] p1_add_3673_comb;
  wire [19:0] p1_concat_3675_comb;
  wire p1_or_3676_comb;
  wire p1_or_3677_comb;
  wire [31:0] p1_add_3716_comb;
  wire [30:0] p1_add_3718_comb;
  wire p1_and_3641_comb;
  wire p1_or_3645_comb;
  wire [31:0] p1_shll_3647_comb;
  wire [31:0] p1_xor_3648_comb;
  wire [31:0] p1_shra_3649_comb;
  wire [31:0] p1_or_3650_comb;
  wire [31:0] p1_sign_ext_3651_comb;
  wire [7:0] p1_array_index_3653_comb;
  wire p1_or_3655_comb;
  wire [31:0] p1_concat_3725_comb;
  wire [31:0] p1_concat_3726_comb;
  wire p1_or_3733_comb;
  wire [3:0] p1_and_3748_comb;
  wire [7:0] p1_array_update_3749_comb[16];
  wire [31:0] p1_add_3751_comb;
  wire [12:0] p1_add_3754_comb;
  wire [8:0] p1_concat_3681_comb;
  wire [8:0] p1_concat_3691_comb;
  wire [10:0] p1_concat_3701_comb;
  wire [5:0] p1_and_3758_comb;
  wire [31:0] p1_add_3759_comb;
  wire [31:0] p1_sel_3760_comb;
  wire [31:0] p1_sel_3761_comb;
  wire [31:0] p1_sel_3762_comb;
  wire [31:0] p1_sel_3763_comb;
  wire [31:0] p1_sel_3764_comb;
  wire [31:0] p1_sel_3765_comb;
  wire [30:0] p1_add_3766_comb;
  wire [7:0] p1_array_update_3774_comb[16];
  wire [31:0] p1_add_3776_comb;
  wire [6:0] p1_concat_3734_comb;
  wire [31:0] p1_sub_3739_comb;
  wire [31:0] p1_add_3740_comb;
  wire [9:0] p1_concat_3781_comb;
  wire [8:0] p1_concat_3790_comb;
  wire [6:0] p1_concat_3800_comb;
  wire [7:0] p1_array_update_3814_comb[16];
  wire [31:0] p1_add_3816_comb;
  wire [7:0] p1_array_update_3817_comb[16];
  wire [3:0] p1_concat_3825_comb;
  wire [7:0] p1_array_update_3826_comb[16];
  wire [7:0] p1_array_update_3827_comb[16];
  wire [7:0] p1_array_update_3828_comb[16];
  wire [4:0] p1_concat_3807_comb;
  wire [31:0] p1_array_update_3808_comb[32];
  wire [31:0] p1_array_update_3809_comb[32];
  wire [31:0] p1_array_update_3810_comb[32];
  wire [31:0] p1_array_update_3811_comb[32];
  wire [31:0] p1_concat_3836_comb;
  wire [7:0] p1_one_hot_sel_3837_comb[16];
  assign p1_bit_slice_3549_comb = p0_ins[31:20];
  assign p1_eq_3551_comb = p0_ins[14:12] == 3'h7;
  assign p1_eq_3552_comb = p0_ins[14:12] == 3'h6;
  assign p1_eq_3553_comb = p0_ins[14:12] == 3'h5;
  assign p1_eq_3554_comb = p0_ins[14:12] == 3'h4;
  assign p1_eq_3555_comb = p0_ins[14:12] == 3'h1;
  assign p1_eq_3556_comb = p0_ins[14:12] == 3'h0;
  assign p1_concat_3557_comb = {20'h0_0000, p1_bit_slice_3549_comb};
  assign p1_array_index_3558_comb = p0_regs[p0_ins[19:15]];
  assign p1_concat_3561_comb = {p1_eq_3551_comb, p1_eq_3552_comb, p1_eq_3553_comb, p1_eq_3553_comb, p1_eq_3554_comb, p1_eq_3555_comb, p1_eq_3556_comb};
  assign p1_add_3564_comb = p1_concat_3557_comb + p1_array_index_3558_comb;
  assign p1_eq_3569_comb = p0_ins[6:0] == 7'h13;
  assign p1_eq_3577_comb = p0_ins[6:0] == 7'h67;
  assign p1_eq_3571_comb = p0_ins[6:0] == 7'h03;
  assign p1_one_hot_3570_comb = {p1_concat_3561_comb[6:0] == 7'h00, p1_concat_3561_comb[6] && p1_concat_3561_comb[5:0] == 6'h00, p1_concat_3561_comb[5] && p1_concat_3561_comb[4:0] == 5'h00, p1_concat_3561_comb[4] && p1_concat_3561_comb[3:0] == 4'h0, p1_concat_3561_comb[3] && p1_concat_3561_comb[2:0] == 3'h0, p1_concat_3561_comb[2] && p1_concat_3561_comb[1:0] == 2'h0, p1_concat_3561_comb[1] && !p1_concat_3561_comb[0], p1_concat_3561_comb[0]};
  assign p1_eq_3572_comb = p0_ins[14:12] == 3'h2;
  assign p1_eq_3594_comb = p0_ins[6:0] == 7'h33;
  assign p1_eq_3595_comb = p0_ins[6:0] == 7'h23;
  assign p1_or_3596_comb = p1_eq_3569_comb | p1_eq_3577_comb | p1_eq_3571_comb;
  assign p1_eq_3597_comb = p0_ins[6:0] == 7'h63;
  assign p1_eq_3598_comb = p0_ins[6:0] == 7'h37;
  assign p1_eq_3599_comb = p0_ins[6:0] == 7'h6f;
  assign p1_add_3587_comb = p1_add_3564_comb[31:1] + 31'h0000_0001;
  assign p1_concat_3612_comb = {p0_ins[31], p0_ins[7], p0_ins[30:25], p0_ins[11:8]};
  assign p1_or_3615_comb = p1_eq_3594_comb | p1_eq_3595_comb | p1_or_3596_comb | p1_eq_3597_comb | p1_eq_3598_comb | p1_eq_3599_comb;
  assign p1_concat_3629_comb = {1'h0, p0_ins[31:25], p0_ins[11:7]};
  assign p1_array_index_3631_comb = p0_regs[p0_ins[24:20]];
  assign p1_concat_3601_comb = {p0_ins[31:25] != 7'h20, p0_ins[31:25] == 7'h20};
  assign p1_and_3602_comb = {7{p1_eq_3569_comb}} & p1_one_hot_3570_comb[6:0];
  assign p1_and_3604_comb = {5{p1_eq_3571_comb}} & {p1_eq_3553_comb, p1_eq_3554_comb, p1_eq_3572_comb, p1_eq_3555_comb, p1_eq_3556_comb};
  assign p1_and_3637_comb = p1_or_3596_comb & ~(p1_eq_3569_comb | p1_eq_3571_comb) & p1_eq_3577_comb & p0_ins[14:12] != 3'h0;
  assign p1_ugt_3667_comb = p0_ins[14:12] > 3'h2;
  assign p1_concat_3668_comb = {20'h0_0000, p0_ins[31:25], p0_ins[11:7]};
  assign p1_add_3670_comb = p1_concat_3629_comb + 13'h0001;
  assign p1_and_3616_comb = {2{p1_eq_3553_comb}} & p1_concat_3601_comb;
  assign p1_array_index_3619_comb = p0_dmem[p1_add_3564_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3564_comb];
  assign p1_add_3620_comb = p1_add_3564_comb + 32'h0000_0001;
  assign p1_array_index_3623_comb = p0_dmem[{p1_add_3587_comb, p1_add_3564_comb[0]} > 32'h0000_000f ? 32'h0000_000f : {p1_add_3587_comb, p1_add_3564_comb[0]}];
  assign p1_add_3624_comb = p1_add_3564_comb + 32'h0000_0003;
  assign p1_add_3626_comb = p0_pc[31:2] + 30'h0000_0001;
  assign p1_add_3673_comb = {{19{p1_concat_3612_comb[11]}}, p1_concat_3612_comb} + p0_pc[31:1];
  assign p1_concat_3675_comb = {p0_ins[31], p0_ins[19:12], p0_ins[20], p0_ins[30:21]};
  assign p1_or_3676_comb = p1_eq_3594_comb | p1_eq_3595_comb | p1_eq_3598_comb | p1_eq_3569_comb | p1_eq_3571_comb;
  assign p1_or_3677_comb = p1_and_3637_comb | ~p1_or_3615_comb;
  assign p1_add_3716_comb = p1_concat_3668_comb + p1_array_index_3631_comb;
  assign p1_add_3718_comb = p1_array_index_3631_comb[31:1] + 31'h0000_0001;
  assign p1_and_3641_comb = p1_eq_3577_comb & p1_eq_3556_comb;
  assign p1_or_3645_comb = p1_and_3602_comb[1] | p1_and_3602_comb[3];
  assign p1_shll_3647_comb = p1_bit_slice_3549_comb >= 12'h020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_bit_slice_3549_comb;
  assign p1_xor_3648_comb = p1_array_index_3558_comb ^ p1_concat_3557_comb;
  assign p1_shra_3649_comb = p1_bit_slice_3549_comb >= 12'h020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_bit_slice_3549_comb);
  assign p1_or_3650_comb = p1_array_index_3558_comb | p1_concat_3557_comb;
  assign p1_sign_ext_3651_comb = {{24{p1_array_index_3619_comb[7]}}, p1_array_index_3619_comb};
  assign p1_array_index_3653_comb = p0_dmem[p1_add_3620_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3620_comb];
  assign p1_or_3655_comb = p1_and_3604_comb[1] | p1_and_3604_comb[4];
  assign p1_concat_3725_comb = {p1_add_3626_comb, p0_pc[1:0]};
  assign p1_concat_3726_comb = {p1_add_3673_comb, p0_pc[0]};
  assign p1_or_3733_comb = p1_or_3676_comb | p1_or_3677_comb;
  assign p1_and_3748_comb = {4{p1_eq_3595_comb}} & {p1_ugt_3667_comb, p1_eq_3556_comb, p1_eq_3555_comb, p1_eq_3572_comb};
  assign p1_array_update_3749_comb[0] = p1_add_3716_comb == 32'h0000_0000 ? p1_array_index_3558_comb[31:24] : p0_dmem[0];
  assign p1_array_update_3749_comb[1] = p1_add_3716_comb == 32'h0000_0001 ? p1_array_index_3558_comb[31:24] : p0_dmem[1];
  assign p1_array_update_3749_comb[2] = p1_add_3716_comb == 32'h0000_0002 ? p1_array_index_3558_comb[31:24] : p0_dmem[2];
  assign p1_array_update_3749_comb[3] = p1_add_3716_comb == 32'h0000_0003 ? p1_array_index_3558_comb[31:24] : p0_dmem[3];
  assign p1_array_update_3749_comb[4] = p1_add_3716_comb == 32'h0000_0004 ? p1_array_index_3558_comb[31:24] : p0_dmem[4];
  assign p1_array_update_3749_comb[5] = p1_add_3716_comb == 32'h0000_0005 ? p1_array_index_3558_comb[31:24] : p0_dmem[5];
  assign p1_array_update_3749_comb[6] = p1_add_3716_comb == 32'h0000_0006 ? p1_array_index_3558_comb[31:24] : p0_dmem[6];
  assign p1_array_update_3749_comb[7] = p1_add_3716_comb == 32'h0000_0007 ? p1_array_index_3558_comb[31:24] : p0_dmem[7];
  assign p1_array_update_3749_comb[8] = p1_add_3716_comb == 32'h0000_0008 ? p1_array_index_3558_comb[31:24] : p0_dmem[8];
  assign p1_array_update_3749_comb[9] = p1_add_3716_comb == 32'h0000_0009 ? p1_array_index_3558_comb[31:24] : p0_dmem[9];
  assign p1_array_update_3749_comb[10] = p1_add_3716_comb == 32'h0000_000a ? p1_array_index_3558_comb[31:24] : p0_dmem[10];
  assign p1_array_update_3749_comb[11] = p1_add_3716_comb == 32'h0000_000b ? p1_array_index_3558_comb[31:24] : p0_dmem[11];
  assign p1_array_update_3749_comb[12] = p1_add_3716_comb == 32'h0000_000c ? p1_array_index_3558_comb[31:24] : p0_dmem[12];
  assign p1_array_update_3749_comb[13] = p1_add_3716_comb == 32'h0000_000d ? p1_array_index_3558_comb[31:24] : p0_dmem[13];
  assign p1_array_update_3749_comb[14] = p1_add_3716_comb == 32'h0000_000e ? p1_array_index_3558_comb[31:24] : p0_dmem[14];
  assign p1_array_update_3749_comb[15] = p1_add_3716_comb == 32'h0000_000f ? p1_array_index_3558_comb[31:24] : p0_dmem[15];
  assign p1_add_3751_comb = {19'h0_0000, p1_add_3670_comb} + p1_array_index_3631_comb;
  assign p1_add_3754_comb = p1_concat_3629_comb + 13'h0003;
  assign p1_concat_3681_comb = {p1_and_3641_comb, p1_and_3604_comb[2:0], p1_and_3602_comb[5:4], p1_and_3602_comb[2], p1_or_3645_comb, p1_and_3602_comb[0]};
  assign p1_concat_3691_comb = {p1_and_3641_comb, p1_and_3604_comb[2], p1_or_3655_comb, p1_and_3604_comb[0], p1_and_3602_comb[5:4], p1_and_3602_comb[2], p1_or_3645_comb, p1_and_3602_comb[0]};
  assign p1_concat_3701_comb = {p1_and_3641_comb, p1_and_3604_comb[3:2], p1_or_3655_comb, p1_and_3604_comb[0], p1_and_3602_comb[6:4], p1_and_3602_comb[2], p1_or_3645_comb, p1_and_3602_comb[0]};
  assign p1_and_3758_comb = {6{p1_eq_3597_comb}} & {p1_eq_3551_comb, p1_eq_3552_comb, p1_eq_3553_comb, p1_eq_3554_comb, p1_eq_3555_comb, p1_eq_3556_comb};
  assign p1_add_3759_comb = {{20{p1_bit_slice_3549_comb[11]}}, p1_bit_slice_3549_comb} + p1_array_index_3558_comb;
  assign p1_sel_3760_comb = p1_array_index_3558_comb == p1_array_index_3631_comb ? p1_concat_3726_comb : p1_concat_3725_comb;
  assign p1_sel_3761_comb = p1_array_index_3558_comb != p1_array_index_3631_comb ? p1_concat_3726_comb : p1_concat_3725_comb;
  assign p1_sel_3762_comb = $signed(p1_array_index_3558_comb) < $signed(p1_array_index_3631_comb) ? p1_concat_3726_comb : p1_concat_3725_comb;
  assign p1_sel_3763_comb = $signed(p1_array_index_3558_comb) >= $signed(p1_array_index_3631_comb) ? p1_concat_3726_comb : p1_concat_3725_comb;
  assign p1_sel_3764_comb = p1_array_index_3558_comb < p1_array_index_3631_comb ? p1_concat_3726_comb : p1_concat_3725_comb;
  assign p1_sel_3765_comb = p1_array_index_3558_comb >= p1_array_index_3631_comb ? p1_concat_3726_comb : p1_concat_3725_comb;
  assign p1_add_3766_comb = {{11{p1_concat_3675_comb[19]}}, p1_concat_3675_comb} + p0_pc[31:1];
  assign p1_array_update_3774_comb[0] = p1_add_3751_comb == 32'h0000_0000 ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[0];
  assign p1_array_update_3774_comb[1] = p1_add_3751_comb == 32'h0000_0001 ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[1];
  assign p1_array_update_3774_comb[2] = p1_add_3751_comb == 32'h0000_0002 ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[2];
  assign p1_array_update_3774_comb[3] = p1_add_3751_comb == 32'h0000_0003 ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[3];
  assign p1_array_update_3774_comb[4] = p1_add_3751_comb == 32'h0000_0004 ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[4];
  assign p1_array_update_3774_comb[5] = p1_add_3751_comb == 32'h0000_0005 ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[5];
  assign p1_array_update_3774_comb[6] = p1_add_3751_comb == 32'h0000_0006 ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[6];
  assign p1_array_update_3774_comb[7] = p1_add_3751_comb == 32'h0000_0007 ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[7];
  assign p1_array_update_3774_comb[8] = p1_add_3751_comb == 32'h0000_0008 ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[8];
  assign p1_array_update_3774_comb[9] = p1_add_3751_comb == 32'h0000_0009 ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[9];
  assign p1_array_update_3774_comb[10] = p1_add_3751_comb == 32'h0000_000a ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[10];
  assign p1_array_update_3774_comb[11] = p1_add_3751_comb == 32'h0000_000b ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[11];
  assign p1_array_update_3774_comb[12] = p1_add_3751_comb == 32'h0000_000c ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[12];
  assign p1_array_update_3774_comb[13] = p1_add_3751_comb == 32'h0000_000d ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[13];
  assign p1_array_update_3774_comb[14] = p1_add_3751_comb == 32'h0000_000e ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[14];
  assign p1_array_update_3774_comb[15] = p1_add_3751_comb == 32'h0000_000f ? p1_array_index_3558_comb[23:16] : p1_array_update_3749_comb[15];
  assign p1_add_3776_comb = p1_concat_3668_comb + {p1_add_3718_comb, p1_array_index_3631_comb[0]};
  assign p1_concat_3734_comb = {p1_and_3616_comb[0], {2{p1_eq_3556_comb}} & p1_concat_3601_comb, p1_eq_3555_comb | p1_and_3616_comb[1], p1_eq_3552_comb, p1_eq_3551_comb, p1_eq_3554_comb};
  assign p1_sub_3739_comb = p1_array_index_3558_comb - p1_array_index_3631_comb;
  assign p1_add_3740_comb = p1_array_index_3631_comb + p1_array_index_3558_comb;
  assign p1_concat_3781_comb = {p1_eq_3599_comb, p1_and_3758_comb, p1_or_3677_comb, p1_and_3641_comb, p1_or_3676_comb};
  assign p1_concat_3790_comb = {p1_eq_3599_comb, p1_and_3758_comb, p1_and_3641_comb, p1_or_3733_comb};
  assign p1_concat_3800_comb = {p1_and_3758_comb, p1_or_3733_comb | p1_eq_3599_comb};
  assign p1_array_update_3814_comb[0] = p1_add_3776_comb == 32'h0000_0000 ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[0];
  assign p1_array_update_3814_comb[1] = p1_add_3776_comb == 32'h0000_0001 ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[1];
  assign p1_array_update_3814_comb[2] = p1_add_3776_comb == 32'h0000_0002 ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[2];
  assign p1_array_update_3814_comb[3] = p1_add_3776_comb == 32'h0000_0003 ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[3];
  assign p1_array_update_3814_comb[4] = p1_add_3776_comb == 32'h0000_0004 ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[4];
  assign p1_array_update_3814_comb[5] = p1_add_3776_comb == 32'h0000_0005 ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[5];
  assign p1_array_update_3814_comb[6] = p1_add_3776_comb == 32'h0000_0006 ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[6];
  assign p1_array_update_3814_comb[7] = p1_add_3776_comb == 32'h0000_0007 ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[7];
  assign p1_array_update_3814_comb[8] = p1_add_3776_comb == 32'h0000_0008 ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[8];
  assign p1_array_update_3814_comb[9] = p1_add_3776_comb == 32'h0000_0009 ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[9];
  assign p1_array_update_3814_comb[10] = p1_add_3776_comb == 32'h0000_000a ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[10];
  assign p1_array_update_3814_comb[11] = p1_add_3776_comb == 32'h0000_000b ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[11];
  assign p1_array_update_3814_comb[12] = p1_add_3776_comb == 32'h0000_000c ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[12];
  assign p1_array_update_3814_comb[13] = p1_add_3776_comb == 32'h0000_000d ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[13];
  assign p1_array_update_3814_comb[14] = p1_add_3776_comb == 32'h0000_000e ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[14];
  assign p1_array_update_3814_comb[15] = p1_add_3776_comb == 32'h0000_000f ? p1_array_index_3558_comb[15:8] : p1_array_update_3774_comb[15];
  assign p1_add_3816_comb = {19'h0_0000, p1_add_3754_comb} + p1_array_index_3631_comb;
  assign p1_array_update_3817_comb[0] = p1_add_3716_comb == 32'h0000_0000 ? p1_array_index_3558_comb[15:8] : p0_dmem[0];
  assign p1_array_update_3817_comb[1] = p1_add_3716_comb == 32'h0000_0001 ? p1_array_index_3558_comb[15:8] : p0_dmem[1];
  assign p1_array_update_3817_comb[2] = p1_add_3716_comb == 32'h0000_0002 ? p1_array_index_3558_comb[15:8] : p0_dmem[2];
  assign p1_array_update_3817_comb[3] = p1_add_3716_comb == 32'h0000_0003 ? p1_array_index_3558_comb[15:8] : p0_dmem[3];
  assign p1_array_update_3817_comb[4] = p1_add_3716_comb == 32'h0000_0004 ? p1_array_index_3558_comb[15:8] : p0_dmem[4];
  assign p1_array_update_3817_comb[5] = p1_add_3716_comb == 32'h0000_0005 ? p1_array_index_3558_comb[15:8] : p0_dmem[5];
  assign p1_array_update_3817_comb[6] = p1_add_3716_comb == 32'h0000_0006 ? p1_array_index_3558_comb[15:8] : p0_dmem[6];
  assign p1_array_update_3817_comb[7] = p1_add_3716_comb == 32'h0000_0007 ? p1_array_index_3558_comb[15:8] : p0_dmem[7];
  assign p1_array_update_3817_comb[8] = p1_add_3716_comb == 32'h0000_0008 ? p1_array_index_3558_comb[15:8] : p0_dmem[8];
  assign p1_array_update_3817_comb[9] = p1_add_3716_comb == 32'h0000_0009 ? p1_array_index_3558_comb[15:8] : p0_dmem[9];
  assign p1_array_update_3817_comb[10] = p1_add_3716_comb == 32'h0000_000a ? p1_array_index_3558_comb[15:8] : p0_dmem[10];
  assign p1_array_update_3817_comb[11] = p1_add_3716_comb == 32'h0000_000b ? p1_array_index_3558_comb[15:8] : p0_dmem[11];
  assign p1_array_update_3817_comb[12] = p1_add_3716_comb == 32'h0000_000c ? p1_array_index_3558_comb[15:8] : p0_dmem[12];
  assign p1_array_update_3817_comb[13] = p1_add_3716_comb == 32'h0000_000d ? p1_array_index_3558_comb[15:8] : p0_dmem[13];
  assign p1_array_update_3817_comb[14] = p1_add_3716_comb == 32'h0000_000e ? p1_array_index_3558_comb[15:8] : p0_dmem[14];
  assign p1_array_update_3817_comb[15] = p1_add_3716_comb == 32'h0000_000f ? p1_array_index_3558_comb[15:8] : p0_dmem[15];
  assign p1_concat_3825_comb = {p1_and_3748_comb[2:0], p0_ins[6:0] != 7'h23 | p1_and_3748_comb[3]};
  assign p1_array_update_3826_comb[0] = p1_add_3816_comb == 32'h0000_0000 ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[0];
  assign p1_array_update_3826_comb[1] = p1_add_3816_comb == 32'h0000_0001 ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[1];
  assign p1_array_update_3826_comb[2] = p1_add_3816_comb == 32'h0000_0002 ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[2];
  assign p1_array_update_3826_comb[3] = p1_add_3816_comb == 32'h0000_0003 ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[3];
  assign p1_array_update_3826_comb[4] = p1_add_3816_comb == 32'h0000_0004 ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[4];
  assign p1_array_update_3826_comb[5] = p1_add_3816_comb == 32'h0000_0005 ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[5];
  assign p1_array_update_3826_comb[6] = p1_add_3816_comb == 32'h0000_0006 ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[6];
  assign p1_array_update_3826_comb[7] = p1_add_3816_comb == 32'h0000_0007 ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[7];
  assign p1_array_update_3826_comb[8] = p1_add_3816_comb == 32'h0000_0008 ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[8];
  assign p1_array_update_3826_comb[9] = p1_add_3816_comb == 32'h0000_0009 ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[9];
  assign p1_array_update_3826_comb[10] = p1_add_3816_comb == 32'h0000_000a ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[10];
  assign p1_array_update_3826_comb[11] = p1_add_3816_comb == 32'h0000_000b ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[11];
  assign p1_array_update_3826_comb[12] = p1_add_3816_comb == 32'h0000_000c ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[12];
  assign p1_array_update_3826_comb[13] = p1_add_3816_comb == 32'h0000_000d ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[13];
  assign p1_array_update_3826_comb[14] = p1_add_3816_comb == 32'h0000_000e ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[14];
  assign p1_array_update_3826_comb[15] = p1_add_3816_comb == 32'h0000_000f ? p1_array_index_3558_comb[7:0] : p1_array_update_3814_comb[15];
  assign p1_array_update_3827_comb[0] = p1_add_3751_comb == 32'h0000_0000 ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[0];
  assign p1_array_update_3827_comb[1] = p1_add_3751_comb == 32'h0000_0001 ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[1];
  assign p1_array_update_3827_comb[2] = p1_add_3751_comb == 32'h0000_0002 ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[2];
  assign p1_array_update_3827_comb[3] = p1_add_3751_comb == 32'h0000_0003 ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[3];
  assign p1_array_update_3827_comb[4] = p1_add_3751_comb == 32'h0000_0004 ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[4];
  assign p1_array_update_3827_comb[5] = p1_add_3751_comb == 32'h0000_0005 ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[5];
  assign p1_array_update_3827_comb[6] = p1_add_3751_comb == 32'h0000_0006 ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[6];
  assign p1_array_update_3827_comb[7] = p1_add_3751_comb == 32'h0000_0007 ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[7];
  assign p1_array_update_3827_comb[8] = p1_add_3751_comb == 32'h0000_0008 ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[8];
  assign p1_array_update_3827_comb[9] = p1_add_3751_comb == 32'h0000_0009 ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[9];
  assign p1_array_update_3827_comb[10] = p1_add_3751_comb == 32'h0000_000a ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[10];
  assign p1_array_update_3827_comb[11] = p1_add_3751_comb == 32'h0000_000b ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[11];
  assign p1_array_update_3827_comb[12] = p1_add_3751_comb == 32'h0000_000c ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[12];
  assign p1_array_update_3827_comb[13] = p1_add_3751_comb == 32'h0000_000d ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[13];
  assign p1_array_update_3827_comb[14] = p1_add_3751_comb == 32'h0000_000e ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[14];
  assign p1_array_update_3827_comb[15] = p1_add_3751_comb == 32'h0000_000f ? p1_array_index_3558_comb[7:0] : p1_array_update_3817_comb[15];
  assign p1_array_update_3828_comb[0] = p1_add_3716_comb == 32'h0000_0000 ? p1_array_index_3558_comb[7:0] : p0_dmem[0];
  assign p1_array_update_3828_comb[1] = p1_add_3716_comb == 32'h0000_0001 ? p1_array_index_3558_comb[7:0] : p0_dmem[1];
  assign p1_array_update_3828_comb[2] = p1_add_3716_comb == 32'h0000_0002 ? p1_array_index_3558_comb[7:0] : p0_dmem[2];
  assign p1_array_update_3828_comb[3] = p1_add_3716_comb == 32'h0000_0003 ? p1_array_index_3558_comb[7:0] : p0_dmem[3];
  assign p1_array_update_3828_comb[4] = p1_add_3716_comb == 32'h0000_0004 ? p1_array_index_3558_comb[7:0] : p0_dmem[4];
  assign p1_array_update_3828_comb[5] = p1_add_3716_comb == 32'h0000_0005 ? p1_array_index_3558_comb[7:0] : p0_dmem[5];
  assign p1_array_update_3828_comb[6] = p1_add_3716_comb == 32'h0000_0006 ? p1_array_index_3558_comb[7:0] : p0_dmem[6];
  assign p1_array_update_3828_comb[7] = p1_add_3716_comb == 32'h0000_0007 ? p1_array_index_3558_comb[7:0] : p0_dmem[7];
  assign p1_array_update_3828_comb[8] = p1_add_3716_comb == 32'h0000_0008 ? p1_array_index_3558_comb[7:0] : p0_dmem[8];
  assign p1_array_update_3828_comb[9] = p1_add_3716_comb == 32'h0000_0009 ? p1_array_index_3558_comb[7:0] : p0_dmem[9];
  assign p1_array_update_3828_comb[10] = p1_add_3716_comb == 32'h0000_000a ? p1_array_index_3558_comb[7:0] : p0_dmem[10];
  assign p1_array_update_3828_comb[11] = p1_add_3716_comb == 32'h0000_000b ? p1_array_index_3558_comb[7:0] : p0_dmem[11];
  assign p1_array_update_3828_comb[12] = p1_add_3716_comb == 32'h0000_000c ? p1_array_index_3558_comb[7:0] : p0_dmem[12];
  assign p1_array_update_3828_comb[13] = p1_add_3716_comb == 32'h0000_000d ? p1_array_index_3558_comb[7:0] : p0_dmem[13];
  assign p1_array_update_3828_comb[14] = p1_add_3716_comb == 32'h0000_000e ? p1_array_index_3558_comb[7:0] : p0_dmem[14];
  assign p1_array_update_3828_comb[15] = p1_add_3716_comb == 32'h0000_000f ? p1_array_index_3558_comb[7:0] : p0_dmem[15];
  assign p1_concat_3807_comb = {p1_eq_3599_comb, p1_eq_3598_comb, p1_or_3596_comb, p1_eq_3595_comb | p1_eq_3597_comb | ~p1_or_3615_comb, p1_eq_3594_comb};
  assign p1_array_update_3808_comb[0] = p0_ins[11:7] == 5'h00 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[0];
  assign p1_array_update_3808_comb[1] = p0_ins[11:7] == 5'h01 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[1];
  assign p1_array_update_3808_comb[2] = p0_ins[11:7] == 5'h02 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[2];
  assign p1_array_update_3808_comb[3] = p0_ins[11:7] == 5'h03 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[3];
  assign p1_array_update_3808_comb[4] = p0_ins[11:7] == 5'h04 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[4];
  assign p1_array_update_3808_comb[5] = p0_ins[11:7] == 5'h05 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[5];
  assign p1_array_update_3808_comb[6] = p0_ins[11:7] == 5'h06 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[6];
  assign p1_array_update_3808_comb[7] = p0_ins[11:7] == 5'h07 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[7];
  assign p1_array_update_3808_comb[8] = p0_ins[11:7] == 5'h08 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[8];
  assign p1_array_update_3808_comb[9] = p0_ins[11:7] == 5'h09 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[9];
  assign p1_array_update_3808_comb[10] = p0_ins[11:7] == 5'h0a ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[10];
  assign p1_array_update_3808_comb[11] = p0_ins[11:7] == 5'h0b ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[11];
  assign p1_array_update_3808_comb[12] = p0_ins[11:7] == 5'h0c ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[12];
  assign p1_array_update_3808_comb[13] = p0_ins[11:7] == 5'h0d ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[13];
  assign p1_array_update_3808_comb[14] = p0_ins[11:7] == 5'h0e ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[14];
  assign p1_array_update_3808_comb[15] = p0_ins[11:7] == 5'h0f ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[15];
  assign p1_array_update_3808_comb[16] = p0_ins[11:7] == 5'h10 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[16];
  assign p1_array_update_3808_comb[17] = p0_ins[11:7] == 5'h11 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[17];
  assign p1_array_update_3808_comb[18] = p0_ins[11:7] == 5'h12 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[18];
  assign p1_array_update_3808_comb[19] = p0_ins[11:7] == 5'h13 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[19];
  assign p1_array_update_3808_comb[20] = p0_ins[11:7] == 5'h14 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[20];
  assign p1_array_update_3808_comb[21] = p0_ins[11:7] == 5'h15 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[21];
  assign p1_array_update_3808_comb[22] = p0_ins[11:7] == 5'h16 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[22];
  assign p1_array_update_3808_comb[23] = p0_ins[11:7] == 5'h17 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[23];
  assign p1_array_update_3808_comb[24] = p0_ins[11:7] == 5'h18 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[24];
  assign p1_array_update_3808_comb[25] = p0_ins[11:7] == 5'h19 ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[25];
  assign p1_array_update_3808_comb[26] = p0_ins[11:7] == 5'h1a ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[26];
  assign p1_array_update_3808_comb[27] = p0_ins[11:7] == 5'h1b ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[27];
  assign p1_array_update_3808_comb[28] = p0_ins[11:7] == 5'h1c ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[28];
  assign p1_array_update_3808_comb[29] = p0_ins[11:7] == 5'h1d ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[29];
  assign p1_array_update_3808_comb[30] = p0_ins[11:7] == 5'h1e ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[30];
  assign p1_array_update_3808_comb[31] = p0_ins[11:7] == 5'h1f ? (p1_array_index_3558_comb ^ p1_array_index_3631_comb) & {32{p1_concat_3734_comb[0]}} | p1_array_index_3558_comb & p1_array_index_3631_comb & {32{p1_concat_3734_comb[1]}} | (p1_array_index_3558_comb | p1_array_index_3631_comb) & {32{p1_concat_3734_comb[2]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? 32'h0000_0000 : p1_array_index_3558_comb << p1_array_index_3631_comb) & {32{p1_concat_3734_comb[3]}} | p1_sub_3739_comb & {32{p1_concat_3734_comb[4]}} | p1_add_3740_comb & {32{p1_concat_3734_comb[5]}} | (p1_array_index_3631_comb >= 32'h0000_0020 ? {32{p1_array_index_3558_comb[31]}} : $unsigned($signed(p1_array_index_3558_comb) >>> p1_array_index_3631_comb)) & {32{p1_concat_3734_comb[6]}} : p0_regs[31];
  assign p1_array_update_3809_comb[0] = p0_ins[11:7] == 5'h00 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[0];
  assign p1_array_update_3809_comb[1] = p0_ins[11:7] == 5'h01 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[1];
  assign p1_array_update_3809_comb[2] = p0_ins[11:7] == 5'h02 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[2];
  assign p1_array_update_3809_comb[3] = p0_ins[11:7] == 5'h03 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[3];
  assign p1_array_update_3809_comb[4] = p0_ins[11:7] == 5'h04 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[4];
  assign p1_array_update_3809_comb[5] = p0_ins[11:7] == 5'h05 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[5];
  assign p1_array_update_3809_comb[6] = p0_ins[11:7] == 5'h06 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[6];
  assign p1_array_update_3809_comb[7] = p0_ins[11:7] == 5'h07 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[7];
  assign p1_array_update_3809_comb[8] = p0_ins[11:7] == 5'h08 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[8];
  assign p1_array_update_3809_comb[9] = p0_ins[11:7] == 5'h09 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[9];
  assign p1_array_update_3809_comb[10] = p0_ins[11:7] == 5'h0a ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[10];
  assign p1_array_update_3809_comb[11] = p0_ins[11:7] == 5'h0b ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[11];
  assign p1_array_update_3809_comb[12] = p0_ins[11:7] == 5'h0c ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[12];
  assign p1_array_update_3809_comb[13] = p0_ins[11:7] == 5'h0d ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[13];
  assign p1_array_update_3809_comb[14] = p0_ins[11:7] == 5'h0e ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[14];
  assign p1_array_update_3809_comb[15] = p0_ins[11:7] == 5'h0f ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[15];
  assign p1_array_update_3809_comb[16] = p0_ins[11:7] == 5'h10 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[16];
  assign p1_array_update_3809_comb[17] = p0_ins[11:7] == 5'h11 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[17];
  assign p1_array_update_3809_comb[18] = p0_ins[11:7] == 5'h12 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[18];
  assign p1_array_update_3809_comb[19] = p0_ins[11:7] == 5'h13 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[19];
  assign p1_array_update_3809_comb[20] = p0_ins[11:7] == 5'h14 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[20];
  assign p1_array_update_3809_comb[21] = p0_ins[11:7] == 5'h15 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[21];
  assign p1_array_update_3809_comb[22] = p0_ins[11:7] == 5'h16 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[22];
  assign p1_array_update_3809_comb[23] = p0_ins[11:7] == 5'h17 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[23];
  assign p1_array_update_3809_comb[24] = p0_ins[11:7] == 5'h18 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[24];
  assign p1_array_update_3809_comb[25] = p0_ins[11:7] == 5'h19 ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[25];
  assign p1_array_update_3809_comb[26] = p0_ins[11:7] == 5'h1a ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[26];
  assign p1_array_update_3809_comb[27] = p0_ins[11:7] == 5'h1b ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[27];
  assign p1_array_update_3809_comb[28] = p0_ins[11:7] == 5'h1c ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[28];
  assign p1_array_update_3809_comb[29] = p0_ins[11:7] == 5'h1d ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[29];
  assign p1_array_update_3809_comb[30] = p0_ins[11:7] == 5'h1e ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[30];
  assign p1_array_update_3809_comb[31] = p0_ins[11:7] == 5'h1f ? {p1_add_3564_comb[31:16] & {16{p1_concat_3681_comb[0]}} | p1_shll_3647_comb[31:16] & {16{p1_concat_3681_comb[1]}} | p1_xor_3648_comb[31:16] & {16{p1_concat_3681_comb[2]}} | p1_shra_3649_comb[31:16] & {16{p1_concat_3681_comb[3]}} | p1_or_3650_comb[31:16] & {16{p1_concat_3681_comb[4]}} | p1_sign_ext_3651_comb[31:16] & {16{p1_concat_3681_comb[5]}} | {16{p1_array_index_3619_comb[7]}} & {16{p1_concat_3681_comb[6]}} | {p1_array_index_3619_comb, p1_array_index_3653_comb} & {16{p1_concat_3681_comb[7]}} | p1_add_3626_comb[29:14] & {16{p1_concat_3681_comb[8]}}, p1_add_3564_comb[15:12] & {4{p1_concat_3691_comb[0]}} | p1_shll_3647_comb[15:12] & {4{p1_concat_3691_comb[1]}} | p1_xor_3648_comb[15:12] & {4{p1_concat_3691_comb[2]}} | p1_shra_3649_comb[15:12] & {4{p1_concat_3691_comb[3]}} | p1_or_3650_comb[15:12] & {4{p1_concat_3691_comb[4]}} | p1_sign_ext_3651_comb[15:12] & {4{p1_concat_3691_comb[5]}} | p1_array_index_3619_comb[7:4] & {4{p1_concat_3691_comb[6]}} | p1_array_index_3623_comb[7:4] & {4{p1_concat_3691_comb[7]}} | p1_add_3626_comb[13:10] & {4{p1_concat_3691_comb[8]}}, p1_add_3564_comb[11:0] & {12{p1_concat_3701_comb[0]}} | p1_shll_3647_comb[11:0] & {12{p1_concat_3701_comb[1]}} | p1_xor_3648_comb[11:0] & {12{p1_concat_3701_comb[2]}} | p1_shra_3649_comb[11:0] & {12{p1_concat_3701_comb[3]}} | p1_or_3650_comb[11:0] & {12{p1_concat_3701_comb[4]}} | p1_array_index_3558_comb[11:0] & p1_bit_slice_3549_comb & {12{p1_concat_3701_comb[5]}} | p1_sign_ext_3651_comb[11:0] & {12{p1_concat_3701_comb[6]}} | {p1_array_index_3619_comb[3:0], p1_array_index_3653_comb} & {12{p1_concat_3701_comb[7]}} | {p1_array_index_3623_comb[3:0], p0_dmem[p1_add_3624_comb > 32'h0000_000f ? 32'h0000_000f : p1_add_3624_comb]} & {12{p1_concat_3701_comb[8]}} | {4'h0, p0_dmem[p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb] > 32'h0000_000f ? 32'h0000_000f : p0_regs[p1_add_3564_comb > 32'h0000_001f ? 32'h0000_001f : p1_add_3564_comb]]} & {12{p1_concat_3701_comb[9]}} | {p1_add_3626_comb[9:0], p0_pc[1:0]} & {12{p1_concat_3701_comb[10]}}} : p0_regs[31];
  assign p1_array_update_3810_comb[0] = p0_ins[11:7] == 5'h00 ? {p0_ins[31:12], 12'h000} : p0_regs[0];
  assign p1_array_update_3810_comb[1] = p0_ins[11:7] == 5'h01 ? {p0_ins[31:12], 12'h000} : p0_regs[1];
  assign p1_array_update_3810_comb[2] = p0_ins[11:7] == 5'h02 ? {p0_ins[31:12], 12'h000} : p0_regs[2];
  assign p1_array_update_3810_comb[3] = p0_ins[11:7] == 5'h03 ? {p0_ins[31:12], 12'h000} : p0_regs[3];
  assign p1_array_update_3810_comb[4] = p0_ins[11:7] == 5'h04 ? {p0_ins[31:12], 12'h000} : p0_regs[4];
  assign p1_array_update_3810_comb[5] = p0_ins[11:7] == 5'h05 ? {p0_ins[31:12], 12'h000} : p0_regs[5];
  assign p1_array_update_3810_comb[6] = p0_ins[11:7] == 5'h06 ? {p0_ins[31:12], 12'h000} : p0_regs[6];
  assign p1_array_update_3810_comb[7] = p0_ins[11:7] == 5'h07 ? {p0_ins[31:12], 12'h000} : p0_regs[7];
  assign p1_array_update_3810_comb[8] = p0_ins[11:7] == 5'h08 ? {p0_ins[31:12], 12'h000} : p0_regs[8];
  assign p1_array_update_3810_comb[9] = p0_ins[11:7] == 5'h09 ? {p0_ins[31:12], 12'h000} : p0_regs[9];
  assign p1_array_update_3810_comb[10] = p0_ins[11:7] == 5'h0a ? {p0_ins[31:12], 12'h000} : p0_regs[10];
  assign p1_array_update_3810_comb[11] = p0_ins[11:7] == 5'h0b ? {p0_ins[31:12], 12'h000} : p0_regs[11];
  assign p1_array_update_3810_comb[12] = p0_ins[11:7] == 5'h0c ? {p0_ins[31:12], 12'h000} : p0_regs[12];
  assign p1_array_update_3810_comb[13] = p0_ins[11:7] == 5'h0d ? {p0_ins[31:12], 12'h000} : p0_regs[13];
  assign p1_array_update_3810_comb[14] = p0_ins[11:7] == 5'h0e ? {p0_ins[31:12], 12'h000} : p0_regs[14];
  assign p1_array_update_3810_comb[15] = p0_ins[11:7] == 5'h0f ? {p0_ins[31:12], 12'h000} : p0_regs[15];
  assign p1_array_update_3810_comb[16] = p0_ins[11:7] == 5'h10 ? {p0_ins[31:12], 12'h000} : p0_regs[16];
  assign p1_array_update_3810_comb[17] = p0_ins[11:7] == 5'h11 ? {p0_ins[31:12], 12'h000} : p0_regs[17];
  assign p1_array_update_3810_comb[18] = p0_ins[11:7] == 5'h12 ? {p0_ins[31:12], 12'h000} : p0_regs[18];
  assign p1_array_update_3810_comb[19] = p0_ins[11:7] == 5'h13 ? {p0_ins[31:12], 12'h000} : p0_regs[19];
  assign p1_array_update_3810_comb[20] = p0_ins[11:7] == 5'h14 ? {p0_ins[31:12], 12'h000} : p0_regs[20];
  assign p1_array_update_3810_comb[21] = p0_ins[11:7] == 5'h15 ? {p0_ins[31:12], 12'h000} : p0_regs[21];
  assign p1_array_update_3810_comb[22] = p0_ins[11:7] == 5'h16 ? {p0_ins[31:12], 12'h000} : p0_regs[22];
  assign p1_array_update_3810_comb[23] = p0_ins[11:7] == 5'h17 ? {p0_ins[31:12], 12'h000} : p0_regs[23];
  assign p1_array_update_3810_comb[24] = p0_ins[11:7] == 5'h18 ? {p0_ins[31:12], 12'h000} : p0_regs[24];
  assign p1_array_update_3810_comb[25] = p0_ins[11:7] == 5'h19 ? {p0_ins[31:12], 12'h000} : p0_regs[25];
  assign p1_array_update_3810_comb[26] = p0_ins[11:7] == 5'h1a ? {p0_ins[31:12], 12'h000} : p0_regs[26];
  assign p1_array_update_3810_comb[27] = p0_ins[11:7] == 5'h1b ? {p0_ins[31:12], 12'h000} : p0_regs[27];
  assign p1_array_update_3810_comb[28] = p0_ins[11:7] == 5'h1c ? {p0_ins[31:12], 12'h000} : p0_regs[28];
  assign p1_array_update_3810_comb[29] = p0_ins[11:7] == 5'h1d ? {p0_ins[31:12], 12'h000} : p0_regs[29];
  assign p1_array_update_3810_comb[30] = p0_ins[11:7] == 5'h1e ? {p0_ins[31:12], 12'h000} : p0_regs[30];
  assign p1_array_update_3810_comb[31] = p0_ins[11:7] == 5'h1f ? {p0_ins[31:12], 12'h000} : p0_regs[31];
  assign p1_array_update_3811_comb[0] = p0_ins[11:7] == 5'h00 ? p1_concat_3725_comb : p0_regs[0];
  assign p1_array_update_3811_comb[1] = p0_ins[11:7] == 5'h01 ? p1_concat_3725_comb : p0_regs[1];
  assign p1_array_update_3811_comb[2] = p0_ins[11:7] == 5'h02 ? p1_concat_3725_comb : p0_regs[2];
  assign p1_array_update_3811_comb[3] = p0_ins[11:7] == 5'h03 ? p1_concat_3725_comb : p0_regs[3];
  assign p1_array_update_3811_comb[4] = p0_ins[11:7] == 5'h04 ? p1_concat_3725_comb : p0_regs[4];
  assign p1_array_update_3811_comb[5] = p0_ins[11:7] == 5'h05 ? p1_concat_3725_comb : p0_regs[5];
  assign p1_array_update_3811_comb[6] = p0_ins[11:7] == 5'h06 ? p1_concat_3725_comb : p0_regs[6];
  assign p1_array_update_3811_comb[7] = p0_ins[11:7] == 5'h07 ? p1_concat_3725_comb : p0_regs[7];
  assign p1_array_update_3811_comb[8] = p0_ins[11:7] == 5'h08 ? p1_concat_3725_comb : p0_regs[8];
  assign p1_array_update_3811_comb[9] = p0_ins[11:7] == 5'h09 ? p1_concat_3725_comb : p0_regs[9];
  assign p1_array_update_3811_comb[10] = p0_ins[11:7] == 5'h0a ? p1_concat_3725_comb : p0_regs[10];
  assign p1_array_update_3811_comb[11] = p0_ins[11:7] == 5'h0b ? p1_concat_3725_comb : p0_regs[11];
  assign p1_array_update_3811_comb[12] = p0_ins[11:7] == 5'h0c ? p1_concat_3725_comb : p0_regs[12];
  assign p1_array_update_3811_comb[13] = p0_ins[11:7] == 5'h0d ? p1_concat_3725_comb : p0_regs[13];
  assign p1_array_update_3811_comb[14] = p0_ins[11:7] == 5'h0e ? p1_concat_3725_comb : p0_regs[14];
  assign p1_array_update_3811_comb[15] = p0_ins[11:7] == 5'h0f ? p1_concat_3725_comb : p0_regs[15];
  assign p1_array_update_3811_comb[16] = p0_ins[11:7] == 5'h10 ? p1_concat_3725_comb : p0_regs[16];
  assign p1_array_update_3811_comb[17] = p0_ins[11:7] == 5'h11 ? p1_concat_3725_comb : p0_regs[17];
  assign p1_array_update_3811_comb[18] = p0_ins[11:7] == 5'h12 ? p1_concat_3725_comb : p0_regs[18];
  assign p1_array_update_3811_comb[19] = p0_ins[11:7] == 5'h13 ? p1_concat_3725_comb : p0_regs[19];
  assign p1_array_update_3811_comb[20] = p0_ins[11:7] == 5'h14 ? p1_concat_3725_comb : p0_regs[20];
  assign p1_array_update_3811_comb[21] = p0_ins[11:7] == 5'h15 ? p1_concat_3725_comb : p0_regs[21];
  assign p1_array_update_3811_comb[22] = p0_ins[11:7] == 5'h16 ? p1_concat_3725_comb : p0_regs[22];
  assign p1_array_update_3811_comb[23] = p0_ins[11:7] == 5'h17 ? p1_concat_3725_comb : p0_regs[23];
  assign p1_array_update_3811_comb[24] = p0_ins[11:7] == 5'h18 ? p1_concat_3725_comb : p0_regs[24];
  assign p1_array_update_3811_comb[25] = p0_ins[11:7] == 5'h19 ? p1_concat_3725_comb : p0_regs[25];
  assign p1_array_update_3811_comb[26] = p0_ins[11:7] == 5'h1a ? p1_concat_3725_comb : p0_regs[26];
  assign p1_array_update_3811_comb[27] = p0_ins[11:7] == 5'h1b ? p1_concat_3725_comb : p0_regs[27];
  assign p1_array_update_3811_comb[28] = p0_ins[11:7] == 5'h1c ? p1_concat_3725_comb : p0_regs[28];
  assign p1_array_update_3811_comb[29] = p0_ins[11:7] == 5'h1d ? p1_concat_3725_comb : p0_regs[29];
  assign p1_array_update_3811_comb[30] = p0_ins[11:7] == 5'h1e ? p1_concat_3725_comb : p0_regs[30];
  assign p1_array_update_3811_comb[31] = p0_ins[11:7] == 5'h1f ? p1_concat_3725_comb : p0_regs[31];
  assign p1_concat_3836_comb = {p1_add_3626_comb & {30{p1_concat_3781_comb[0]}} | p1_add_3759_comb[31:2] & {30{p1_concat_3781_comb[1]}} | p0_pc[31:2] & {30{p1_concat_3781_comb[2]}} | p1_sel_3760_comb[31:2] & {30{p1_concat_3781_comb[3]}} | p1_sel_3761_comb[31:2] & {30{p1_concat_3781_comb[4]}} | p1_sel_3762_comb[31:2] & {30{p1_concat_3781_comb[5]}} | p1_sel_3763_comb[31:2] & {30{p1_concat_3781_comb[6]}} | p1_sel_3764_comb[31:2] & {30{p1_concat_3781_comb[7]}} | p1_sel_3765_comb[31:2] & {30{p1_concat_3781_comb[8]}} | p1_add_3766_comb[30:1] & {30{p1_concat_3781_comb[9]}}, p0_pc[1] & p1_concat_3790_comb[0] | p1_add_3759_comb[1] & p1_concat_3790_comb[1] | p1_sel_3760_comb[1] & p1_concat_3790_comb[2] | p1_sel_3761_comb[1] & p1_concat_3790_comb[3] | p1_sel_3762_comb[1] & p1_concat_3790_comb[4] | p1_sel_3763_comb[1] & p1_concat_3790_comb[5] | p1_sel_3764_comb[1] & p1_concat_3790_comb[6] | p1_sel_3765_comb[1] & p1_concat_3790_comb[7] | p1_add_3766_comb[0] & p1_concat_3790_comb[8], p0_pc[0] & p1_concat_3800_comb[0] | p1_sel_3760_comb[0] & p1_concat_3800_comb[1] | p1_sel_3761_comb[0] & p1_concat_3800_comb[2] | p1_sel_3762_comb[0] & p1_concat_3800_comb[3] | p1_sel_3763_comb[0] & p1_concat_3800_comb[4] | p1_sel_3764_comb[0] & p1_concat_3800_comb[5] | p1_sel_3765_comb[0] & p1_concat_3800_comb[6]};
  assign p1_one_hot_sel_3837_comb[0] = p0_dmem[0] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[0] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[0] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[0] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[1] = p0_dmem[1] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[1] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[1] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[1] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[2] = p0_dmem[2] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[2] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[2] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[2] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[3] = p0_dmem[3] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[3] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[3] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[3] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[4] = p0_dmem[4] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[4] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[4] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[4] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[5] = p0_dmem[5] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[5] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[5] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[5] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[6] = p0_dmem[6] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[6] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[6] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[6] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[7] = p0_dmem[7] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[7] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[7] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[7] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[8] = p0_dmem[8] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[8] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[8] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[8] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[9] = p0_dmem[9] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[9] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[9] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[9] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[10] = p0_dmem[10] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[10] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[10] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[10] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[11] = p0_dmem[11] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[11] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[11] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[11] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[12] = p0_dmem[12] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[12] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[12] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[12] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[13] = p0_dmem[13] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[13] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[13] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[13] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[14] = p0_dmem[14] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[14] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[14] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[14] & {8{p1_concat_3825_comb[3]}};
  assign p1_one_hot_sel_3837_comb[15] = p0_dmem[15] & {8{p1_concat_3825_comb[0]}} | p1_array_update_3826_comb[15] & {8{p1_concat_3825_comb[1]}} | p1_array_update_3827_comb[15] & {8{p1_concat_3825_comb[2]}} | p1_array_update_3828_comb[15] & {8{p1_concat_3825_comb[3]}};

  // Registers for pipe stage 1:
  reg [31:0] p1_regs[32];
  reg [4:0] p1_concat_3807;
  reg [31:0] p1_array_update_3808[32];
  reg [31:0] p1_array_update_3809[32];
  reg [31:0] p1_array_update_3810[32];
  reg [31:0] p1_array_update_3811[32];
  reg [31:0] p1_concat_3836;
  reg [7:0] p1_one_hot_sel_3837[16];
  always_ff @ (posedge clk) begin
    p1_regs <= p0_regs;
    p1_concat_3807 <= p1_concat_3807_comb;
    p1_array_update_3808 <= p1_array_update_3808_comb;
    p1_array_update_3809 <= p1_array_update_3809_comb;
    p1_array_update_3810 <= p1_array_update_3810_comb;
    p1_array_update_3811 <= p1_array_update_3811_comb;
    p1_concat_3836 <= p1_concat_3836_comb;
    p1_one_hot_sel_3837 <= p1_one_hot_sel_3837_comb;
  end

  // ===== Pipe stage 2:
  wire [31:0] p2_one_hot_sel_3861_comb[32];
  assign p2_one_hot_sel_3861_comb[0] = p1_array_update_3808[0] & {32{p1_concat_3807[0]}} | p1_regs[0] & {32{p1_concat_3807[1]}} | p1_array_update_3809[0] & {32{p1_concat_3807[2]}} | p1_array_update_3810[0] & {32{p1_concat_3807[3]}} | p1_array_update_3811[0] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[1] = p1_array_update_3808[1] & {32{p1_concat_3807[0]}} | p1_regs[1] & {32{p1_concat_3807[1]}} | p1_array_update_3809[1] & {32{p1_concat_3807[2]}} | p1_array_update_3810[1] & {32{p1_concat_3807[3]}} | p1_array_update_3811[1] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[2] = p1_array_update_3808[2] & {32{p1_concat_3807[0]}} | p1_regs[2] & {32{p1_concat_3807[1]}} | p1_array_update_3809[2] & {32{p1_concat_3807[2]}} | p1_array_update_3810[2] & {32{p1_concat_3807[3]}} | p1_array_update_3811[2] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[3] = p1_array_update_3808[3] & {32{p1_concat_3807[0]}} | p1_regs[3] & {32{p1_concat_3807[1]}} | p1_array_update_3809[3] & {32{p1_concat_3807[2]}} | p1_array_update_3810[3] & {32{p1_concat_3807[3]}} | p1_array_update_3811[3] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[4] = p1_array_update_3808[4] & {32{p1_concat_3807[0]}} | p1_regs[4] & {32{p1_concat_3807[1]}} | p1_array_update_3809[4] & {32{p1_concat_3807[2]}} | p1_array_update_3810[4] & {32{p1_concat_3807[3]}} | p1_array_update_3811[4] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[5] = p1_array_update_3808[5] & {32{p1_concat_3807[0]}} | p1_regs[5] & {32{p1_concat_3807[1]}} | p1_array_update_3809[5] & {32{p1_concat_3807[2]}} | p1_array_update_3810[5] & {32{p1_concat_3807[3]}} | p1_array_update_3811[5] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[6] = p1_array_update_3808[6] & {32{p1_concat_3807[0]}} | p1_regs[6] & {32{p1_concat_3807[1]}} | p1_array_update_3809[6] & {32{p1_concat_3807[2]}} | p1_array_update_3810[6] & {32{p1_concat_3807[3]}} | p1_array_update_3811[6] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[7] = p1_array_update_3808[7] & {32{p1_concat_3807[0]}} | p1_regs[7] & {32{p1_concat_3807[1]}} | p1_array_update_3809[7] & {32{p1_concat_3807[2]}} | p1_array_update_3810[7] & {32{p1_concat_3807[3]}} | p1_array_update_3811[7] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[8] = p1_array_update_3808[8] & {32{p1_concat_3807[0]}} | p1_regs[8] & {32{p1_concat_3807[1]}} | p1_array_update_3809[8] & {32{p1_concat_3807[2]}} | p1_array_update_3810[8] & {32{p1_concat_3807[3]}} | p1_array_update_3811[8] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[9] = p1_array_update_3808[9] & {32{p1_concat_3807[0]}} | p1_regs[9] & {32{p1_concat_3807[1]}} | p1_array_update_3809[9] & {32{p1_concat_3807[2]}} | p1_array_update_3810[9] & {32{p1_concat_3807[3]}} | p1_array_update_3811[9] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[10] = p1_array_update_3808[10] & {32{p1_concat_3807[0]}} | p1_regs[10] & {32{p1_concat_3807[1]}} | p1_array_update_3809[10] & {32{p1_concat_3807[2]}} | p1_array_update_3810[10] & {32{p1_concat_3807[3]}} | p1_array_update_3811[10] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[11] = p1_array_update_3808[11] & {32{p1_concat_3807[0]}} | p1_regs[11] & {32{p1_concat_3807[1]}} | p1_array_update_3809[11] & {32{p1_concat_3807[2]}} | p1_array_update_3810[11] & {32{p1_concat_3807[3]}} | p1_array_update_3811[11] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[12] = p1_array_update_3808[12] & {32{p1_concat_3807[0]}} | p1_regs[12] & {32{p1_concat_3807[1]}} | p1_array_update_3809[12] & {32{p1_concat_3807[2]}} | p1_array_update_3810[12] & {32{p1_concat_3807[3]}} | p1_array_update_3811[12] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[13] = p1_array_update_3808[13] & {32{p1_concat_3807[0]}} | p1_regs[13] & {32{p1_concat_3807[1]}} | p1_array_update_3809[13] & {32{p1_concat_3807[2]}} | p1_array_update_3810[13] & {32{p1_concat_3807[3]}} | p1_array_update_3811[13] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[14] = p1_array_update_3808[14] & {32{p1_concat_3807[0]}} | p1_regs[14] & {32{p1_concat_3807[1]}} | p1_array_update_3809[14] & {32{p1_concat_3807[2]}} | p1_array_update_3810[14] & {32{p1_concat_3807[3]}} | p1_array_update_3811[14] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[15] = p1_array_update_3808[15] & {32{p1_concat_3807[0]}} | p1_regs[15] & {32{p1_concat_3807[1]}} | p1_array_update_3809[15] & {32{p1_concat_3807[2]}} | p1_array_update_3810[15] & {32{p1_concat_3807[3]}} | p1_array_update_3811[15] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[16] = p1_array_update_3808[16] & {32{p1_concat_3807[0]}} | p1_regs[16] & {32{p1_concat_3807[1]}} | p1_array_update_3809[16] & {32{p1_concat_3807[2]}} | p1_array_update_3810[16] & {32{p1_concat_3807[3]}} | p1_array_update_3811[16] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[17] = p1_array_update_3808[17] & {32{p1_concat_3807[0]}} | p1_regs[17] & {32{p1_concat_3807[1]}} | p1_array_update_3809[17] & {32{p1_concat_3807[2]}} | p1_array_update_3810[17] & {32{p1_concat_3807[3]}} | p1_array_update_3811[17] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[18] = p1_array_update_3808[18] & {32{p1_concat_3807[0]}} | p1_regs[18] & {32{p1_concat_3807[1]}} | p1_array_update_3809[18] & {32{p1_concat_3807[2]}} | p1_array_update_3810[18] & {32{p1_concat_3807[3]}} | p1_array_update_3811[18] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[19] = p1_array_update_3808[19] & {32{p1_concat_3807[0]}} | p1_regs[19] & {32{p1_concat_3807[1]}} | p1_array_update_3809[19] & {32{p1_concat_3807[2]}} | p1_array_update_3810[19] & {32{p1_concat_3807[3]}} | p1_array_update_3811[19] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[20] = p1_array_update_3808[20] & {32{p1_concat_3807[0]}} | p1_regs[20] & {32{p1_concat_3807[1]}} | p1_array_update_3809[20] & {32{p1_concat_3807[2]}} | p1_array_update_3810[20] & {32{p1_concat_3807[3]}} | p1_array_update_3811[20] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[21] = p1_array_update_3808[21] & {32{p1_concat_3807[0]}} | p1_regs[21] & {32{p1_concat_3807[1]}} | p1_array_update_3809[21] & {32{p1_concat_3807[2]}} | p1_array_update_3810[21] & {32{p1_concat_3807[3]}} | p1_array_update_3811[21] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[22] = p1_array_update_3808[22] & {32{p1_concat_3807[0]}} | p1_regs[22] & {32{p1_concat_3807[1]}} | p1_array_update_3809[22] & {32{p1_concat_3807[2]}} | p1_array_update_3810[22] & {32{p1_concat_3807[3]}} | p1_array_update_3811[22] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[23] = p1_array_update_3808[23] & {32{p1_concat_3807[0]}} | p1_regs[23] & {32{p1_concat_3807[1]}} | p1_array_update_3809[23] & {32{p1_concat_3807[2]}} | p1_array_update_3810[23] & {32{p1_concat_3807[3]}} | p1_array_update_3811[23] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[24] = p1_array_update_3808[24] & {32{p1_concat_3807[0]}} | p1_regs[24] & {32{p1_concat_3807[1]}} | p1_array_update_3809[24] & {32{p1_concat_3807[2]}} | p1_array_update_3810[24] & {32{p1_concat_3807[3]}} | p1_array_update_3811[24] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[25] = p1_array_update_3808[25] & {32{p1_concat_3807[0]}} | p1_regs[25] & {32{p1_concat_3807[1]}} | p1_array_update_3809[25] & {32{p1_concat_3807[2]}} | p1_array_update_3810[25] & {32{p1_concat_3807[3]}} | p1_array_update_3811[25] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[26] = p1_array_update_3808[26] & {32{p1_concat_3807[0]}} | p1_regs[26] & {32{p1_concat_3807[1]}} | p1_array_update_3809[26] & {32{p1_concat_3807[2]}} | p1_array_update_3810[26] & {32{p1_concat_3807[3]}} | p1_array_update_3811[26] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[27] = p1_array_update_3808[27] & {32{p1_concat_3807[0]}} | p1_regs[27] & {32{p1_concat_3807[1]}} | p1_array_update_3809[27] & {32{p1_concat_3807[2]}} | p1_array_update_3810[27] & {32{p1_concat_3807[3]}} | p1_array_update_3811[27] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[28] = p1_array_update_3808[28] & {32{p1_concat_3807[0]}} | p1_regs[28] & {32{p1_concat_3807[1]}} | p1_array_update_3809[28] & {32{p1_concat_3807[2]}} | p1_array_update_3810[28] & {32{p1_concat_3807[3]}} | p1_array_update_3811[28] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[29] = p1_array_update_3808[29] & {32{p1_concat_3807[0]}} | p1_regs[29] & {32{p1_concat_3807[1]}} | p1_array_update_3809[29] & {32{p1_concat_3807[2]}} | p1_array_update_3810[29] & {32{p1_concat_3807[3]}} | p1_array_update_3811[29] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[30] = p1_array_update_3808[30] & {32{p1_concat_3807[0]}} | p1_regs[30] & {32{p1_concat_3807[1]}} | p1_array_update_3809[30] & {32{p1_concat_3807[2]}} | p1_array_update_3810[30] & {32{p1_concat_3807[3]}} | p1_array_update_3811[30] & {32{p1_concat_3807[4]}};
  assign p2_one_hot_sel_3861_comb[31] = p1_array_update_3808[31] & {32{p1_concat_3807[0]}} | p1_regs[31] & {32{p1_concat_3807[1]}} | p1_array_update_3809[31] & {32{p1_concat_3807[2]}} | p1_array_update_3810[31] & {32{p1_concat_3807[3]}} | p1_array_update_3811[31] & {32{p1_concat_3807[4]}};

  // Registers for pipe stage 2:
  reg [31:0] p2_one_hot_sel_3861[32];
  reg [31:0] p2_concat_3836;
  reg [7:0] p2_one_hot_sel_3837[16];
  always_ff @ (posedge clk) begin
    p2_one_hot_sel_3861 <= p2_one_hot_sel_3861_comb;
    p2_concat_3836 <= p1_concat_3836;
    p2_one_hot_sel_3837 <= p1_one_hot_sel_3837;
  end

  // ===== Pipe stage 3:
  wire [31:0] p3_array_update_3870_comb[32];
  wire [1183:0] p3_tuple_3871_comb;
  assign p3_array_update_3870_comb[0] = 32'h0000_0000;
  assign p3_array_update_3870_comb[1] = p2_one_hot_sel_3861[1];
  assign p3_array_update_3870_comb[2] = p2_one_hot_sel_3861[2];
  assign p3_array_update_3870_comb[3] = p2_one_hot_sel_3861[3];
  assign p3_array_update_3870_comb[4] = p2_one_hot_sel_3861[4];
  assign p3_array_update_3870_comb[5] = p2_one_hot_sel_3861[5];
  assign p3_array_update_3870_comb[6] = p2_one_hot_sel_3861[6];
  assign p3_array_update_3870_comb[7] = p2_one_hot_sel_3861[7];
  assign p3_array_update_3870_comb[8] = p2_one_hot_sel_3861[8];
  assign p3_array_update_3870_comb[9] = p2_one_hot_sel_3861[9];
  assign p3_array_update_3870_comb[10] = p2_one_hot_sel_3861[10];
  assign p3_array_update_3870_comb[11] = p2_one_hot_sel_3861[11];
  assign p3_array_update_3870_comb[12] = p2_one_hot_sel_3861[12];
  assign p3_array_update_3870_comb[13] = p2_one_hot_sel_3861[13];
  assign p3_array_update_3870_comb[14] = p2_one_hot_sel_3861[14];
  assign p3_array_update_3870_comb[15] = p2_one_hot_sel_3861[15];
  assign p3_array_update_3870_comb[16] = p2_one_hot_sel_3861[16];
  assign p3_array_update_3870_comb[17] = p2_one_hot_sel_3861[17];
  assign p3_array_update_3870_comb[18] = p2_one_hot_sel_3861[18];
  assign p3_array_update_3870_comb[19] = p2_one_hot_sel_3861[19];
  assign p3_array_update_3870_comb[20] = p2_one_hot_sel_3861[20];
  assign p3_array_update_3870_comb[21] = p2_one_hot_sel_3861[21];
  assign p3_array_update_3870_comb[22] = p2_one_hot_sel_3861[22];
  assign p3_array_update_3870_comb[23] = p2_one_hot_sel_3861[23];
  assign p3_array_update_3870_comb[24] = p2_one_hot_sel_3861[24];
  assign p3_array_update_3870_comb[25] = p2_one_hot_sel_3861[25];
  assign p3_array_update_3870_comb[26] = p2_one_hot_sel_3861[26];
  assign p3_array_update_3870_comb[27] = p2_one_hot_sel_3861[27];
  assign p3_array_update_3870_comb[28] = p2_one_hot_sel_3861[28];
  assign p3_array_update_3870_comb[29] = p2_one_hot_sel_3861[29];
  assign p3_array_update_3870_comb[30] = p2_one_hot_sel_3861[30];
  assign p3_array_update_3870_comb[31] = p2_one_hot_sel_3861[31];
  assign p3_tuple_3871_comb = {p2_concat_3836, {p3_array_update_3870_comb[31], p3_array_update_3870_comb[30], p3_array_update_3870_comb[29], p3_array_update_3870_comb[28], p3_array_update_3870_comb[27], p3_array_update_3870_comb[26], p3_array_update_3870_comb[25], p3_array_update_3870_comb[24], p3_array_update_3870_comb[23], p3_array_update_3870_comb[22], p3_array_update_3870_comb[21], p3_array_update_3870_comb[20], p3_array_update_3870_comb[19], p3_array_update_3870_comb[18], p3_array_update_3870_comb[17], p3_array_update_3870_comb[16], p3_array_update_3870_comb[15], p3_array_update_3870_comb[14], p3_array_update_3870_comb[13], p3_array_update_3870_comb[12], p3_array_update_3870_comb[11], p3_array_update_3870_comb[10], p3_array_update_3870_comb[9], p3_array_update_3870_comb[8], p3_array_update_3870_comb[7], p3_array_update_3870_comb[6], p3_array_update_3870_comb[5], p3_array_update_3870_comb[4], p3_array_update_3870_comb[3], p3_array_update_3870_comb[2], p3_array_update_3870_comb[1], p3_array_update_3870_comb[0]}, {p2_one_hot_sel_3837[15], p2_one_hot_sel_3837[14], p2_one_hot_sel_3837[13], p2_one_hot_sel_3837[12], p2_one_hot_sel_3837[11], p2_one_hot_sel_3837[10], p2_one_hot_sel_3837[9], p2_one_hot_sel_3837[8], p2_one_hot_sel_3837[7], p2_one_hot_sel_3837[6], p2_one_hot_sel_3837[5], p2_one_hot_sel_3837[4], p2_one_hot_sel_3837[3], p2_one_hot_sel_3837[2], p2_one_hot_sel_3837[1], p2_one_hot_sel_3837[0]}};

  // Registers for pipe stage 3:
  reg [1183:0] p3_tuple_3871;
  always_ff @ (posedge clk) begin
    p3_tuple_3871 <= p3_tuple_3871_comb;
  end
  __riscv_simple__run_instruction_13___itok__riscv_simple__run_instruction_unsupported_func3: assert property (@(posedge clk) disable iff ($isunknown(p1_or_3615_comb)) p1_or_3615_comb) else $fatal(0, "Assertion failure via fail! @ xls/examples/riscv_simple.x:535:17-535:56");
  unmatched_func3: assert property (@(posedge clk) disable iff ($isunknown(~(p1_eq_3594_comb & ~(p1_eq_3554_comb | p1_eq_3551_comb | p1_eq_3552_comb | p1_eq_3555_comb | p1_eq_3556_comb | p1_eq_3553_comb)))) ~(p1_eq_3594_comb & ~(p1_eq_3554_comb | p1_eq_3551_comb | p1_eq_3552_comb | p1_eq_3555_comb | p1_eq_3556_comb | p1_eq_3553_comb))) else $fatal(0, "Assertion failure via fail! @ xls/examples/riscv_simple.x:372:18-372:44");
  unsupported_funct3: assert property (@(posedge clk) disable iff ($isunknown(~(p1_eq_3595_comb & p1_ugt_3667_comb))) ~(p1_eq_3595_comb & p1_ugt_3667_comb)) else $fatal(0, "Assertion failure via fail! @ xls/examples/riscv_simple.x:468:21-468:49");
  unmatched_I_ARITH_func3: assert property (@(posedge clk) disable iff ($isunknown(~(p1_or_3596_comb & p1_eq_3569_comb & ~(p1_eq_3554_comb | p1_eq_3551_comb | p1_eq_3552_comb | p1_eq_3555_comb | p1_eq_3556_comb | p1_eq_3553_comb)))) ~(p1_or_3596_comb & p1_eq_3569_comb & ~(p1_eq_3554_comb | p1_eq_3551_comb | p1_eq_3552_comb | p1_eq_3555_comb | p1_eq_3556_comb | p1_eq_3553_comb))) else $fatal(0, "Assertion failure via fail! @ xls/examples/riscv_simple.x:396:25-396:59");
  unmatched_I_LD_func3: assert property (@(posedge clk) disable iff ($isunknown(~(p1_or_3596_comb & p0_ins[6:0] != 7'h13 & p1_eq_3571_comb & ~(p1_eq_3556_comb | p1_eq_3555_comb | p1_eq_3572_comb | p1_eq_3554_comb | p1_eq_3553_comb)))) ~(p1_or_3596_comb & p0_ins[6:0] != 7'h13 & p1_eq_3571_comb & ~(p1_eq_3556_comb | p1_eq_3555_comb | p1_eq_3572_comb | p1_eq_3554_comb | p1_eq_3553_comb))) else $fatal(0, "Assertion failure via fail! @ xls/examples/riscv_simple.x:413:25-413:56");
  unmatched_I_JALR_funct3: assert property (@(posedge clk) disable iff ($isunknown(~p1_and_3637_comb)) ~p1_and_3637_comb) else $fatal(0, "Assertion failure via fail! @ xls/examples/riscv_simple.x:423:26-423:66");
  __riscv_simple__run_instruction_13___itok__riscv_simple__run_instruction___itok__riscv_simple__run_instruction_10___itok__riscv_simple__run_b_instruction_unsupported_func3: assert property (@(posedge clk) disable iff ($isunknown(~(p1_eq_3597_comb & ~(p1_eq_3554_comb | p1_eq_3551_comb | p1_eq_3552_comb | p1_eq_3555_comb | p1_eq_3556_comb | p1_eq_3553_comb)))) ~(p1_eq_3597_comb & ~(p1_eq_3554_comb | p1_eq_3551_comb | p1_eq_3552_comb | p1_eq_3555_comb | p1_eq_3556_comb | p1_eq_3553_comb))) else $fatal(0, "Assertion failure via fail! @ xls/examples/riscv_simple.x:512:19-512:47");
  assign out = p3_tuple_3871;
endmodule
