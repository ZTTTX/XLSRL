module xls_test(
  input wire clk,
  input wire [2047:0] f,
  output wire [2047:0] out
);
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_11b (input reg [31:0] lhs, input reg [10:0] rhs);
    begin
      umul32b_32b_x_11b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_12b (input reg [31:0] lhs, input reg [11:0] rhs);
    begin
      umul32b_32b_x_12b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_10b (input reg [31:0] lhs, input reg [9:0] rhs);
    begin
      umul32b_32b_x_10b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  // lint_off MULTIPLY
  function automatic [31:0] umul32b_32b_x_8b (input reg [31:0] lhs, input reg [7:0] rhs);
    begin
      umul32b_32b_x_8b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [31:0] f_unflattened[64];
  assign f_unflattened[0] = f[31:0];
  assign f_unflattened[1] = f[63:32];
  assign f_unflattened[2] = f[95:64];
  assign f_unflattened[3] = f[127:96];
  assign f_unflattened[4] = f[159:128];
  assign f_unflattened[5] = f[191:160];
  assign f_unflattened[6] = f[223:192];
  assign f_unflattened[7] = f[255:224];
  assign f_unflattened[8] = f[287:256];
  assign f_unflattened[9] = f[319:288];
  assign f_unflattened[10] = f[351:320];
  assign f_unflattened[11] = f[383:352];
  assign f_unflattened[12] = f[415:384];
  assign f_unflattened[13] = f[447:416];
  assign f_unflattened[14] = f[479:448];
  assign f_unflattened[15] = f[511:480];
  assign f_unflattened[16] = f[543:512];
  assign f_unflattened[17] = f[575:544];
  assign f_unflattened[18] = f[607:576];
  assign f_unflattened[19] = f[639:608];
  assign f_unflattened[20] = f[671:640];
  assign f_unflattened[21] = f[703:672];
  assign f_unflattened[22] = f[735:704];
  assign f_unflattened[23] = f[767:736];
  assign f_unflattened[24] = f[799:768];
  assign f_unflattened[25] = f[831:800];
  assign f_unflattened[26] = f[863:832];
  assign f_unflattened[27] = f[895:864];
  assign f_unflattened[28] = f[927:896];
  assign f_unflattened[29] = f[959:928];
  assign f_unflattened[30] = f[991:960];
  assign f_unflattened[31] = f[1023:992];
  assign f_unflattened[32] = f[1055:1024];
  assign f_unflattened[33] = f[1087:1056];
  assign f_unflattened[34] = f[1119:1088];
  assign f_unflattened[35] = f[1151:1120];
  assign f_unflattened[36] = f[1183:1152];
  assign f_unflattened[37] = f[1215:1184];
  assign f_unflattened[38] = f[1247:1216];
  assign f_unflattened[39] = f[1279:1248];
  assign f_unflattened[40] = f[1311:1280];
  assign f_unflattened[41] = f[1343:1312];
  assign f_unflattened[42] = f[1375:1344];
  assign f_unflattened[43] = f[1407:1376];
  assign f_unflattened[44] = f[1439:1408];
  assign f_unflattened[45] = f[1471:1440];
  assign f_unflattened[46] = f[1503:1472];
  assign f_unflattened[47] = f[1535:1504];
  assign f_unflattened[48] = f[1567:1536];
  assign f_unflattened[49] = f[1599:1568];
  assign f_unflattened[50] = f[1631:1600];
  assign f_unflattened[51] = f[1663:1632];
  assign f_unflattened[52] = f[1695:1664];
  assign f_unflattened[53] = f[1727:1696];
  assign f_unflattened[54] = f[1759:1728];
  assign f_unflattened[55] = f[1791:1760];
  assign f_unflattened[56] = f[1823:1792];
  assign f_unflattened[57] = f[1855:1824];
  assign f_unflattened[58] = f[1887:1856];
  assign f_unflattened[59] = f[1919:1888];
  assign f_unflattened[60] = f[1951:1920];
  assign f_unflattened[61] = f[1983:1952];
  assign f_unflattened[62] = f[2015:1984];
  assign f_unflattened[63] = f[2047:2016];

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_f[64];
  always_ff @ (posedge clk) begin
    p0_f <= f_unflattened;
  end

  // ===== Pipe stage 1:
  wire [31:0] p1_array_index_33119_comb;
  wire [31:0] p1_array_index_33120_comb;
  wire [31:0] p1_array_index_33121_comb;
  wire [31:0] p1_array_index_33122_comb;
  wire [31:0] p1_array_index_33163_comb;
  wire [31:0] p1_array_index_33164_comb;
  wire [31:0] p1_array_index_33165_comb;
  wire [31:0] p1_array_index_33166_comb;
  wire [31:0] p1_array_index_33399_comb;
  wire [31:0] p1_array_index_33400_comb;
  wire [31:0] p1_array_index_33401_comb;
  wire [31:0] p1_array_index_33402_comb;
  wire [31:0] p1_array_index_32895_comb;
  wire [31:0] p1_array_index_32896_comb;
  wire [31:0] p1_array_index_32897_comb;
  wire [31:0] p1_array_index_32898_comb;
  wire [31:0] p1_array_index_32913_comb;
  wire [31:0] p1_array_index_32914_comb;
  wire [31:0] p1_array_index_32915_comb;
  wire [31:0] p1_array_index_32916_comb;
  wire [31:0] p1_array_index_33025_comb;
  wire [31:0] p1_array_index_33026_comb;
  wire [31:0] p1_array_index_33027_comb;
  wire [31:0] p1_array_index_33028_comb;
  wire [31:0] p1_add_33144_comb;
  wire [31:0] p1_add_33147_comb;
  wire [31:0] p1_add_33188_comb;
  wire [31:0] p1_add_33191_comb;
  wire [31:0] p1_add_33468_comb;
  wire [31:0] p1_add_33471_comb;
  wire [31:0] p1_add_32906_comb;
  wire [31:0] p1_add_32911_comb;
  wire [31:0] p1_add_32928_comb;
  wire [31:0] p1_add_32933_comb;
  wire [31:0] p1_add_33052_comb;
  wire [31:0] p1_add_33057_comb;
  wire [31:0] p1_array_index_32917_comb;
  wire [31:0] p1_array_index_32918_comb;
  wire [31:0] p1_array_index_32921_comb;
  wire [31:0] p1_array_index_32922_comb;
  wire [31:0] p1_umul_33167_comb;
  wire [31:0] p1_umul_33168_comb;
  wire [31:0] p1_umul_33169_comb;
  wire [31:0] p1_umul_33170_comb;
  wire [31:0] p1_array_index_32945_comb;
  wire [31:0] p1_array_index_32946_comb;
  wire [31:0] p1_array_index_32949_comb;
  wire [31:0] p1_array_index_32950_comb;
  wire [31:0] p1_umul_33217_comb;
  wire [31:0] p1_umul_33218_comb;
  wire [31:0] p1_umul_33219_comb;
  wire [31:0] p1_umul_33220_comb;
  wire [31:0] p1_array_index_33073_comb;
  wire [31:0] p1_array_index_33074_comb;
  wire [31:0] p1_array_index_33077_comb;
  wire [31:0] p1_array_index_33078_comb;
  wire [31:0] p1_umul_33519_comb;
  wire [31:0] p1_umul_33520_comb;
  wire [31:0] p1_umul_33521_comb;
  wire [31:0] p1_umul_33522_comb;
  wire [31:0] p1_umul_32919_comb;
  wire [31:0] p1_umul_32920_comb;
  wire [31:0] p1_umul_32923_comb;
  wire [31:0] p1_umul_32924_comb;
  wire [31:0] p1_umul_32947_comb;
  wire [31:0] p1_umul_32948_comb;
  wire [31:0] p1_umul_32951_comb;
  wire [31:0] p1_umul_32952_comb;
  wire [31:0] p1_umul_33075_comb;
  wire [31:0] p1_umul_33076_comb;
  wire [31:0] p1_umul_33079_comb;
  wire [31:0] p1_umul_33080_comb;
  wire [31:0] p1_add_32935_comb;
  wire [31:0] p1_add_32940_comb;
  wire [31:0] p1_add_32965_comb;
  wire [31:0] p1_add_32970_comb;
  wire [31:0] p1_add_33101_comb;
  wire [31:0] p1_add_33106_comb;
  wire [31:0] p1_umul_32953_comb;
  wire [20:0] p1_bit_slice_33213_comb;
  wire [20:0] p1_bit_slice_33214_comb;
  wire [31:0] p1_umul_32979_comb;
  wire [31:0] p1_umul_32954_comb;
  wire [31:0] p1_umul_32959_comb;
  wire [20:0] p1_bit_slice_33215_comb;
  wire [20:0] p1_bit_slice_33216_comb;
  wire [31:0] p1_umul_32984_comb;
  wire [31:0] p1_umul_32960_comb;
  wire [31:0] p1_umul_32977_comb;
  wire [26:0] p1_add_33221_comb;
  wire [31:0] p1_umul_32982_comb;
  wire [26:0] p1_add_33222_comb;
  wire [31:0] p1_umul_32985_comb;
  wire [20:0] p1_bit_slice_33293_comb;
  wire [20:0] p1_bit_slice_33294_comb;
  wire [31:0] p1_umul_33013_comb;
  wire [31:0] p1_umul_32986_comb;
  wire [31:0] p1_umul_32991_comb;
  wire [20:0] p1_bit_slice_33295_comb;
  wire [20:0] p1_bit_slice_33296_comb;
  wire [31:0] p1_umul_33018_comb;
  wire [31:0] p1_umul_32992_comb;
  wire [31:0] p1_umul_33011_comb;
  wire [26:0] p1_add_33321_comb;
  wire [31:0] p1_umul_33016_comb;
  wire [26:0] p1_add_33322_comb;
  wire [31:0] p1_umul_33123_comb;
  wire [20:0] p1_bit_slice_33593_comb;
  wire [20:0] p1_bit_slice_33594_comb;
  wire [31:0] p1_umul_33153_comb;
  wire [31:0] p1_umul_33124_comb;
  wire [31:0] p1_umul_33129_comb;
  wire [20:0] p1_bit_slice_33595_comb;
  wire [20:0] p1_bit_slice_33596_comb;
  wire [31:0] p1_umul_33158_comb;
  wire [31:0] p1_umul_33130_comb;
  wire [31:0] p1_umul_33151_comb;
  wire [26:0] p1_add_33597_comb;
  wire [31:0] p1_umul_33156_comb;
  wire [26:0] p1_add_33598_comb;
  wire [29:0] p1_add_32956_comb;
  wire [29:0] p1_add_32962_comb;
  wire [29:0] p1_add_32988_comb;
  wire [29:0] p1_add_32994_comb;
  wire [29:0] p1_add_33126_comb;
  wire [29:0] p1_add_33132_comb;
  wire [20:0] p1_add_33248_comb;
  wire [20:0] p1_add_33254_comb;
  wire [20:0] p1_add_33354_comb;
  wire [20:0] p1_add_33360_comb;
  wire [20:0] p1_add_33610_comb;
  wire [20:0] p1_add_33616_comb;
  wire [31:0] p1_concat_32978_comb;
  wire [31:0] p1_concat_32983_comb;
  wire [31:0] p1_concat_33012_comb;
  wire [31:0] p1_concat_33017_comb;
  wire [31:0] p1_concat_33152_comb;
  wire [31:0] p1_concat_33157_comb;
  wire [24:0] p1_add_33297_comb;
  wire [20:0] p1_add_33299_comb;
  wire [30:0] p1_add_33301_comb;
  wire [24:0] p1_add_33303_comb;
  wire [20:0] p1_add_33305_comb;
  wire [30:0] p1_add_33307_comb;
  wire [24:0] p1_add_33309_comb;
  wire [20:0] p1_add_33311_comb;
  wire [28:0] p1_add_33313_comb;
  wire [24:0] p1_add_33315_comb;
  wire [20:0] p1_add_33317_comb;
  wire [28:0] p1_add_33319_comb;
  wire [24:0] p1_add_33323_comb;
  wire [20:0] p1_add_33325_comb;
  wire [28:0] p1_add_33327_comb;
  wire [24:0] p1_add_33329_comb;
  wire [20:0] p1_add_33331_comb;
  wire [28:0] p1_add_33333_comb;
  wire [24:0] p1_add_33411_comb;
  wire [20:0] p1_add_33413_comb;
  wire [30:0] p1_add_33415_comb;
  wire [24:0] p1_add_33417_comb;
  wire [20:0] p1_add_33419_comb;
  wire [30:0] p1_add_33421_comb;
  wire [24:0] p1_add_33433_comb;
  wire [20:0] p1_add_33435_comb;
  wire [28:0] p1_add_33437_comb;
  wire [24:0] p1_add_33439_comb;
  wire [20:0] p1_add_33441_comb;
  wire [28:0] p1_add_33443_comb;
  wire [24:0] p1_add_33449_comb;
  wire [20:0] p1_add_33451_comb;
  wire [28:0] p1_add_33453_comb;
  wire [24:0] p1_add_33455_comb;
  wire [20:0] p1_add_33457_comb;
  wire [28:0] p1_add_33459_comb;
  wire [24:0] p1_add_33645_comb;
  wire [20:0] p1_add_33647_comb;
  wire [30:0] p1_add_33649_comb;
  wire [24:0] p1_add_33651_comb;
  wire [20:0] p1_add_33653_comb;
  wire [30:0] p1_add_33655_comb;
  wire [24:0] p1_add_33657_comb;
  wire [20:0] p1_add_33659_comb;
  wire [28:0] p1_add_33661_comb;
  wire [24:0] p1_add_33663_comb;
  wire [20:0] p1_add_33665_comb;
  wire [28:0] p1_add_33667_comb;
  wire [24:0] p1_add_33669_comb;
  wire [20:0] p1_add_33671_comb;
  wire [28:0] p1_add_33673_comb;
  wire [24:0] p1_add_33675_comb;
  wire [20:0] p1_add_33677_comb;
  wire [28:0] p1_add_33679_comb;
  wire [28:0] p1_add_32997_comb;
  wire [31:0] p1_add_32999_comb;
  wire [31:0] p1_add_33000_comb;
  wire [28:0] p1_add_33001_comb;
  wire [31:0] p1_add_33003_comb;
  wire [31:0] p1_add_33004_comb;
  wire [28:0] p1_add_33033_comb;
  wire [31:0] p1_add_33035_comb;
  wire [31:0] p1_add_33036_comb;
  wire [28:0] p1_add_33037_comb;
  wire [31:0] p1_add_33039_comb;
  wire [31:0] p1_add_33040_comb;
  wire [28:0] p1_add_33171_comb;
  wire [31:0] p1_add_33173_comb;
  wire [31:0] p1_add_33174_comb;
  wire [28:0] p1_add_33175_comb;
  wire [31:0] p1_add_33177_comb;
  wire [31:0] p1_add_33178_comb;
  wire [31:0] p1_sub_33345_comb;
  wire [31:0] p1_sub_33348_comb;
  wire [29:0] p1_concat_33366_comb;
  wire [29:0] p1_concat_33370_comb;
  wire [31:0] p1_sub_33473_comb;
  wire [31:0] p1_sub_33476_comb;
  wire [29:0] p1_concat_33486_comb;
  wire [29:0] p1_concat_33490_comb;
  wire [31:0] p1_sub_33683_comb;
  wire [31:0] p1_sub_33686_comb;
  wire [29:0] p1_concat_33692_comb;
  wire [29:0] p1_concat_33696_comb;
  wire [31:0] p1_add_33405_comb;
  wire [24:0] p1_add_33406_comb;
  wire [31:0] p1_add_33408_comb;
  wire [24:0] p1_add_33409_comb;
  wire [28:0] p1_add_33423_comb;
  wire [29:0] p1_add_33425_comb;
  wire [28:0] p1_add_33428_comb;
  wire [29:0] p1_add_33430_comb;
  wire [30:0] p1_add_33445_comb;
  wire [29:0] p1_add_33446_comb;
  wire [30:0] p1_add_33447_comb;
  wire [29:0] p1_add_33448_comb;
  wire [29:0] p1_add_33461_comb;
  wire [29:0] p1_add_33463_comb;
  wire [29:0] p1_add_33464_comb;
  wire [29:0] p1_add_33466_comb;
  wire [31:0] p1_add_33523_comb;
  wire [24:0] p1_add_33524_comb;
  wire [31:0] p1_add_33526_comb;
  wire [24:0] p1_add_33527_comb;
  wire [28:0] p1_add_33531_comb;
  wire [29:0] p1_add_33533_comb;
  wire [28:0] p1_add_33536_comb;
  wire [29:0] p1_add_33538_comb;
  wire [30:0] p1_add_33543_comb;
  wire [29:0] p1_add_33544_comb;
  wire [30:0] p1_add_33545_comb;
  wire [29:0] p1_add_33546_comb;
  wire [29:0] p1_add_33549_comb;
  wire [29:0] p1_add_33551_comb;
  wire [29:0] p1_add_33552_comb;
  wire [29:0] p1_add_33554_comb;
  wire [31:0] p1_add_33713_comb;
  wire [24:0] p1_add_33714_comb;
  wire [31:0] p1_add_33716_comb;
  wire [24:0] p1_add_33717_comb;
  wire [28:0] p1_add_33719_comb;
  wire [29:0] p1_add_33721_comb;
  wire [28:0] p1_add_33724_comb;
  wire [29:0] p1_add_33726_comb;
  wire [30:0] p1_add_33729_comb;
  wire [29:0] p1_add_33730_comb;
  wire [30:0] p1_add_33731_comb;
  wire [29:0] p1_add_33732_comb;
  wire [29:0] p1_add_33733_comb;
  wire [29:0] p1_add_33735_comb;
  wire [29:0] p1_add_33736_comb;
  wire [29:0] p1_add_33738_comb;
  wire [28:0] p1_add_33029_comb;
  wire [28:0] p1_add_33031_comb;
  wire [30:0] p1_add_33041_comb;
  wire [28:0] p1_add_33043_comb;
  wire [30:0] p1_add_33045_comb;
  wire [28:0] p1_add_33047_comb;
  wire [28:0] p1_add_33081_comb;
  wire [28:0] p1_add_33083_comb;
  wire [30:0] p1_add_33087_comb;
  wire [28:0] p1_add_33089_comb;
  wire [30:0] p1_add_33091_comb;
  wire [28:0] p1_add_33093_comb;
  wire [28:0] p1_add_33223_comb;
  wire [28:0] p1_add_33225_comb;
  wire [30:0] p1_add_33227_comb;
  wire [28:0] p1_add_33229_comb;
  wire [30:0] p1_add_33231_comb;
  wire [28:0] p1_add_33233_comb;
  wire [31:0] p1_add_33059_comb;
  wire [31:0] p1_add_33061_comb;
  wire [31:0] p1_add_33111_comb;
  wire [31:0] p1_add_33113_comb;
  wire [31:0] p1_add_33277_comb;
  wire [31:0] p1_add_33279_comb;
  wire [29:0] p1_add_33529_comb;
  wire [29:0] p1_add_33530_comb;
  wire [31:0] p1_sub_33541_comb;
  wire [31:0] p1_sub_33542_comb;
  wire [31:0] p1_sub_33547_comb;
  wire [31:0] p1_sub_33548_comb;
  wire [31:0] p1_sub_33555_comb;
  wire [31:0] p1_sub_33556_comb;
  wire [29:0] p1_add_33599_comb;
  wire [29:0] p1_add_33600_comb;
  wire [31:0] p1_sub_33601_comb;
  wire [31:0] p1_sub_33602_comb;
  wire [31:0] p1_sub_33603_comb;
  wire [31:0] p1_sub_33604_comb;
  wire [31:0] p1_sub_33605_comb;
  wire [31:0] p1_sub_33606_comb;
  wire [29:0] p1_add_33759_comb;
  wire [29:0] p1_add_33760_comb;
  wire [31:0] p1_sub_33761_comb;
  wire [31:0] p1_sub_33762_comb;
  wire [31:0] p1_sub_33763_comb;
  wire [31:0] p1_sub_33764_comb;
  wire [31:0] p1_sub_33765_comb;
  wire [31:0] p1_sub_33766_comb;
  wire [31:0] p1_sub_33085_comb;
  wire [31:0] p1_sub_33086_comb;
  wire [31:0] p1_sub_33095_comb;
  wire [31:0] p1_sub_33096_comb;
  wire [31:0] p1_sub_33135_comb;
  wire [31:0] p1_sub_33136_comb;
  wire [31:0] p1_sub_33137_comb;
  wire [31:0] p1_sub_33138_comb;
  wire [31:0] p1_array_index_33203_comb;
  wire [31:0] p1_array_index_33204_comb;
  wire [31:0] p1_array_index_33237_comb;
  wire [31:0] p1_array_index_33238_comb;
  wire [31:0] p1_array_index_33285_comb;
  wire [31:0] p1_array_index_33286_comb;
  wire [31:0] p1_sub_33335_comb;
  wire [31:0] p1_sub_33336_comb;
  wire [31:0] p1_sub_33337_comb;
  wire [31:0] p1_sub_33338_comb;
  wire [31:0] p1_array_index_33343_comb;
  wire [31:0] p1_array_index_33344_comb;
  wire [23:0] p1_bit_slice_33571_comb;
  wire [23:0] p1_bit_slice_33572_comb;
  wire [23:0] p1_bit_slice_33577_comb;
  wire [23:0] p1_bit_slice_33578_comb;
  wire [23:0] p1_bit_slice_33583_comb;
  wire [23:0] p1_bit_slice_33584_comb;
  wire [23:0] p1_bit_slice_33589_comb;
  wire [23:0] p1_bit_slice_33590_comb;
  wire [23:0] p1_bit_slice_33635_comb;
  wire [23:0] p1_bit_slice_33636_comb;
  wire [23:0] p1_bit_slice_33637_comb;
  wire [23:0] p1_bit_slice_33638_comb;
  wire [23:0] p1_bit_slice_33639_comb;
  wire [23:0] p1_bit_slice_33640_comb;
  wire [23:0] p1_bit_slice_33641_comb;
  wire [23:0] p1_bit_slice_33642_comb;
  wire [31:0] p1_array_index_33709_comb;
  wire [31:0] p1_array_index_33710_comb;
  wire [31:0] p1_array_index_33739_comb;
  wire [31:0] p1_array_index_33740_comb;
  wire [23:0] p1_bit_slice_33771_comb;
  wire [23:0] p1_bit_slice_33772_comb;
  wire [23:0] p1_bit_slice_33773_comb;
  wire [23:0] p1_bit_slice_33774_comb;
  wire [23:0] p1_bit_slice_33775_comb;
  wire [23:0] p1_bit_slice_33776_comb;
  wire [23:0] p1_bit_slice_33777_comb;
  wire [23:0] p1_bit_slice_33778_comb;
  wire [20:0] p1_bit_slice_33779_comb;
  wire [20:0] p1_bit_slice_33780_comb;
  wire [20:0] p1_bit_slice_33783_comb;
  wire [20:0] p1_bit_slice_33784_comb;
  wire [31:0] p1_umul_33207_comb;
  wire [31:0] p1_umul_33208_comb;
  wire [31:0] p1_umul_33291_comb;
  wire [31:0] p1_umul_33292_comb;
  wire [31:0] p1_umul_33591_comb;
  wire [31:0] p1_umul_33592_comb;
  assign p1_array_index_33119_comb = p0_f[6'h0a];
  assign p1_array_index_33120_comb = p0_f[6'h0e];
  assign p1_array_index_33121_comb = p0_f[6'h3a];
  assign p1_array_index_33122_comb = p0_f[6'h3e];
  assign p1_array_index_33163_comb = p0_f[6'h2a];
  assign p1_array_index_33164_comb = p0_f[6'h2e];
  assign p1_array_index_33165_comb = p0_f[6'h1a];
  assign p1_array_index_33166_comb = p0_f[6'h1e];
  assign p1_array_index_33399_comb = p0_f[6'h12];
  assign p1_array_index_33400_comb = p0_f[6'h16];
  assign p1_array_index_33401_comb = p0_f[6'h32];
  assign p1_array_index_33402_comb = p0_f[6'h36];
  assign p1_array_index_32895_comb = p0_f[6'h09];
  assign p1_array_index_32896_comb = p0_f[6'h0f];
  assign p1_array_index_32897_comb = p0_f[6'h39];
  assign p1_array_index_32898_comb = p0_f[6'h3f];
  assign p1_array_index_32913_comb = p0_f[6'h29];
  assign p1_array_index_32914_comb = p0_f[6'h2f];
  assign p1_array_index_32915_comb = p0_f[6'h19];
  assign p1_array_index_32916_comb = p0_f[6'h1f];
  assign p1_array_index_33025_comb = p0_f[6'h11];
  assign p1_array_index_33026_comb = p0_f[6'h17];
  assign p1_array_index_33027_comb = p0_f[6'h31];
  assign p1_array_index_33028_comb = p0_f[6'h37];
  assign p1_add_33144_comb = p1_array_index_33119_comb + p1_array_index_33120_comb;
  assign p1_add_33147_comb = p1_array_index_33121_comb + p1_array_index_33122_comb;
  assign p1_add_33188_comb = p1_array_index_33163_comb + p1_array_index_33164_comb;
  assign p1_add_33191_comb = p1_array_index_33165_comb + p1_array_index_33166_comb;
  assign p1_add_33468_comb = p1_array_index_33399_comb + p1_array_index_33400_comb;
  assign p1_add_33471_comb = p1_array_index_33401_comb + p1_array_index_33402_comb;
  assign p1_add_32906_comb = p1_array_index_32895_comb + p1_array_index_32896_comb;
  assign p1_add_32911_comb = p1_array_index_32897_comb + p1_array_index_32898_comb;
  assign p1_add_32928_comb = p1_array_index_32913_comb + p1_array_index_32914_comb;
  assign p1_add_32933_comb = p1_array_index_32915_comb + p1_array_index_32916_comb;
  assign p1_add_33052_comb = p1_array_index_33025_comb + p1_array_index_33026_comb;
  assign p1_add_33057_comb = p1_array_index_33027_comb + p1_array_index_33028_comb;
  assign p1_array_index_32917_comb = p0_f[6'h0d];
  assign p1_array_index_32918_comb = p0_f[6'h0b];
  assign p1_array_index_32921_comb = p0_f[6'h3d];
  assign p1_array_index_32922_comb = p0_f[6'h3b];
  assign p1_umul_33167_comb = umul32b_32b_x_11b(p1_array_index_33119_comb, 11'h620);
  assign p1_umul_33168_comb = umul32b_32b_x_11b(p1_add_33144_comb, 11'h454);
  assign p1_umul_33169_comb = umul32b_32b_x_11b(p1_array_index_33121_comb, 11'h620);
  assign p1_umul_33170_comb = umul32b_32b_x_11b(p1_add_33147_comb, 11'h454);
  assign p1_array_index_32945_comb = p0_f[6'h2d];
  assign p1_array_index_32946_comb = p0_f[6'h2b];
  assign p1_array_index_32949_comb = p0_f[6'h1d];
  assign p1_array_index_32950_comb = p0_f[6'h1b];
  assign p1_umul_33217_comb = umul32b_32b_x_11b(p1_array_index_33163_comb, 11'h620);
  assign p1_umul_33218_comb = umul32b_32b_x_11b(p1_add_33188_comb, 11'h454);
  assign p1_umul_33219_comb = umul32b_32b_x_11b(p1_array_index_33165_comb, 11'h620);
  assign p1_umul_33220_comb = umul32b_32b_x_11b(p1_add_33191_comb, 11'h454);
  assign p1_array_index_33073_comb = p0_f[6'h15];
  assign p1_array_index_33074_comb = p0_f[6'h13];
  assign p1_array_index_33077_comb = p0_f[6'h35];
  assign p1_array_index_33078_comb = p0_f[6'h33];
  assign p1_umul_33519_comb = umul32b_32b_x_11b(p1_array_index_33399_comb, 11'h620);
  assign p1_umul_33520_comb = umul32b_32b_x_11b(p1_add_33468_comb, 11'h454);
  assign p1_umul_33521_comb = umul32b_32b_x_11b(p1_array_index_33401_comb, 11'h620);
  assign p1_umul_33522_comb = umul32b_32b_x_11b(p1_add_33471_comb, 11'h454);
  assign p1_umul_32919_comb = umul32b_32b_x_12b(p1_array_index_32895_comb, 12'h8e4);
  assign p1_umul_32920_comb = umul32b_32b_x_10b(p1_add_32906_comb, 10'h235);
  assign p1_umul_32923_comb = umul32b_32b_x_12b(p1_array_index_32897_comb, 12'h8e4);
  assign p1_umul_32924_comb = umul32b_32b_x_10b(p1_add_32911_comb, 10'h235);
  assign p1_umul_32947_comb = umul32b_32b_x_12b(p1_array_index_32913_comb, 12'h8e4);
  assign p1_umul_32948_comb = umul32b_32b_x_10b(p1_add_32928_comb, 10'h235);
  assign p1_umul_32951_comb = umul32b_32b_x_12b(p1_array_index_32915_comb, 12'h8e4);
  assign p1_umul_32952_comb = umul32b_32b_x_10b(p1_add_32933_comb, 10'h235);
  assign p1_umul_33075_comb = umul32b_32b_x_12b(p1_array_index_33025_comb, 12'h8e4);
  assign p1_umul_33076_comb = umul32b_32b_x_10b(p1_add_33052_comb, 10'h235);
  assign p1_umul_33079_comb = umul32b_32b_x_12b(p1_array_index_33027_comb, 12'h8e4);
  assign p1_umul_33080_comb = umul32b_32b_x_10b(p1_add_33057_comb, 10'h235);
  assign p1_add_32935_comb = p1_array_index_32917_comb + p1_array_index_32918_comb;
  assign p1_add_32940_comb = p1_array_index_32921_comb + p1_array_index_32922_comb;
  assign p1_add_32965_comb = p1_array_index_32945_comb + p1_array_index_32946_comb;
  assign p1_add_32970_comb = p1_array_index_32949_comb + p1_array_index_32950_comb;
  assign p1_add_33101_comb = p1_array_index_33073_comb + p1_array_index_33074_comb;
  assign p1_add_33106_comb = p1_array_index_33077_comb + p1_array_index_33078_comb;
  assign p1_umul_32953_comb = umul32b_32b_x_12b(p1_add_32935_comb, 12'h968);
  assign p1_bit_slice_33213_comb = p0_f[6'h0c][20:0];
  assign p1_bit_slice_33214_comb = p0_f[6'h08][20:0];
  assign p1_umul_32979_comb = umul32b_32b_x_12b(p1_array_index_32918_comb, 12'hfb1);
  assign p1_umul_32954_comb = umul32b_32b_x_12b(p1_array_index_32896_comb, 12'hd4e);
  assign p1_umul_32959_comb = umul32b_32b_x_12b(p1_add_32940_comb, 12'h968);
  assign p1_bit_slice_33215_comb = p0_f[6'h3c][20:0];
  assign p1_bit_slice_33216_comb = p0_f[6'h38][20:0];
  assign p1_umul_32984_comb = umul32b_32b_x_12b(p1_array_index_32922_comb, 12'hfb1);
  assign p1_umul_32960_comb = umul32b_32b_x_12b(p1_array_index_32898_comb, 12'hd4e);
  assign p1_umul_32977_comb = umul32b_32b_x_10b(p1_array_index_32917_comb, 10'h31f);
  assign p1_add_33221_comb = p1_umul_33167_comb[31:5] + p1_umul_33168_comb[31:5];
  assign p1_umul_32982_comb = umul32b_32b_x_10b(p1_array_index_32921_comb, 10'h31f);
  assign p1_add_33222_comb = p1_umul_33169_comb[31:5] + p1_umul_33170_comb[31:5];
  assign p1_umul_32985_comb = umul32b_32b_x_12b(p1_add_32965_comb, 12'h968);
  assign p1_bit_slice_33293_comb = p0_f[6'h2c][20:0];
  assign p1_bit_slice_33294_comb = p0_f[6'h28][20:0];
  assign p1_umul_33013_comb = umul32b_32b_x_12b(p1_array_index_32946_comb, 12'hfb1);
  assign p1_umul_32986_comb = umul32b_32b_x_12b(p1_array_index_32914_comb, 12'hd4e);
  assign p1_umul_32991_comb = umul32b_32b_x_12b(p1_add_32970_comb, 12'h968);
  assign p1_bit_slice_33295_comb = p0_f[6'h1c][20:0];
  assign p1_bit_slice_33296_comb = p0_f[6'h18][20:0];
  assign p1_umul_33018_comb = umul32b_32b_x_12b(p1_array_index_32950_comb, 12'hfb1);
  assign p1_umul_32992_comb = umul32b_32b_x_12b(p1_array_index_32916_comb, 12'hd4e);
  assign p1_umul_33011_comb = umul32b_32b_x_10b(p1_array_index_32945_comb, 10'h31f);
  assign p1_add_33321_comb = p1_umul_33217_comb[31:5] + p1_umul_33218_comb[31:5];
  assign p1_umul_33016_comb = umul32b_32b_x_10b(p1_array_index_32949_comb, 10'h31f);
  assign p1_add_33322_comb = p1_umul_33219_comb[31:5] + p1_umul_33220_comb[31:5];
  assign p1_umul_33123_comb = umul32b_32b_x_12b(p1_add_33101_comb, 12'h968);
  assign p1_bit_slice_33593_comb = p0_f[6'h14][20:0];
  assign p1_bit_slice_33594_comb = p0_f[6'h10][20:0];
  assign p1_umul_33153_comb = umul32b_32b_x_12b(p1_array_index_33074_comb, 12'hfb1);
  assign p1_umul_33124_comb = umul32b_32b_x_12b(p1_array_index_33026_comb, 12'hd4e);
  assign p1_umul_33129_comb = umul32b_32b_x_12b(p1_add_33106_comb, 12'h968);
  assign p1_bit_slice_33595_comb = p0_f[6'h34][20:0];
  assign p1_bit_slice_33596_comb = p0_f[6'h30][20:0];
  assign p1_umul_33158_comb = umul32b_32b_x_12b(p1_array_index_33078_comb, 12'hfb1);
  assign p1_umul_33130_comb = umul32b_32b_x_12b(p1_array_index_33028_comb, 12'hd4e);
  assign p1_umul_33151_comb = umul32b_32b_x_10b(p1_array_index_33073_comb, 10'h31f);
  assign p1_add_33597_comb = p1_umul_33519_comb[31:5] + p1_umul_33520_comb[31:5];
  assign p1_umul_33156_comb = umul32b_32b_x_10b(p1_array_index_33077_comb, 10'h31f);
  assign p1_add_33598_comb = p1_umul_33521_comb[31:5] + p1_umul_33522_comb[31:5];
  assign p1_add_32956_comb = p1_umul_32919_comb[31:2] + p1_umul_32920_comb[31:2];
  assign p1_add_32962_comb = p1_umul_32923_comb[31:2] + p1_umul_32924_comb[31:2];
  assign p1_add_32988_comb = p1_umul_32947_comb[31:2] + p1_umul_32948_comb[31:2];
  assign p1_add_32994_comb = p1_umul_32951_comb[31:2] + p1_umul_32952_comb[31:2];
  assign p1_add_33126_comb = p1_umul_33075_comb[31:2] + p1_umul_33076_comb[31:2];
  assign p1_add_33132_comb = p1_umul_33079_comb[31:2] + p1_umul_33080_comb[31:2];
  assign p1_add_33248_comb = p1_bit_slice_33213_comb + p1_bit_slice_33214_comb;
  assign p1_add_33254_comb = p1_bit_slice_33215_comb + p1_bit_slice_33216_comb;
  assign p1_add_33354_comb = p1_bit_slice_33293_comb + p1_bit_slice_33294_comb;
  assign p1_add_33360_comb = p1_bit_slice_33295_comb + p1_bit_slice_33296_comb;
  assign p1_add_33610_comb = p1_bit_slice_33593_comb + p1_bit_slice_33594_comb;
  assign p1_add_33616_comb = p1_bit_slice_33595_comb + p1_bit_slice_33596_comb;
  assign p1_concat_32978_comb = {p1_add_32956_comb, p1_umul_32920_comb[1:0]};
  assign p1_concat_32983_comb = {p1_add_32962_comb, p1_umul_32924_comb[1:0]};
  assign p1_concat_33012_comb = {p1_add_32988_comb, p1_umul_32948_comb[1:0]};
  assign p1_concat_33017_comb = {p1_add_32994_comb, p1_umul_32952_comb[1:0]};
  assign p1_concat_33152_comb = {p1_add_33126_comb, p1_umul_33076_comb[1:0]};
  assign p1_concat_33157_comb = {p1_add_33132_comb, p1_umul_33080_comb[1:0]};
  assign p1_add_33297_comb = p1_umul_32953_comb[31:7] + 25'h000_0001;
  assign p1_add_33299_comb = p1_umul_32920_comb[31:11] + p1_add_33248_comb;
  assign p1_add_33301_comb = p1_umul_32979_comb[31:1] + p1_umul_32954_comb[31:1];
  assign p1_add_33303_comb = p1_umul_32959_comb[31:7] + 25'h000_0001;
  assign p1_add_33305_comb = p1_umul_32924_comb[31:11] + p1_add_33254_comb;
  assign p1_add_33307_comb = p1_umul_32984_comb[31:1] + p1_umul_32960_comb[31:1];
  assign p1_add_33309_comb = p1_umul_32979_comb[31:7] + 25'h000_0001;
  assign p1_add_33311_comb = p1_umul_32954_comb[31:11] + p1_add_33248_comb;
  assign p1_add_33313_comb = p1_umul_32953_comb[31:3] + p1_umul_32920_comb[31:3];
  assign p1_add_33315_comb = p1_umul_32984_comb[31:7] + 25'h000_0001;
  assign p1_add_33317_comb = p1_umul_32960_comb[31:11] + p1_add_33254_comb;
  assign p1_add_33319_comb = p1_umul_32959_comb[31:3] + p1_umul_32924_comb[31:3];
  assign p1_add_33323_comb = p1_umul_32977_comb[31:7] + 25'h000_0001;
  assign p1_add_33325_comb = p1_add_33221_comb[26:6] + p1_add_33248_comb;
  assign p1_add_33327_comb = p1_umul_32953_comb[31:3] + p1_umul_32919_comb[31:3];
  assign p1_add_33329_comb = p1_umul_32982_comb[31:7] + 25'h000_0001;
  assign p1_add_33331_comb = p1_add_33222_comb[26:6] + p1_add_33254_comb;
  assign p1_add_33333_comb = p1_umul_32959_comb[31:3] + p1_umul_32923_comb[31:3];
  assign p1_add_33411_comb = p1_umul_32985_comb[31:7] + 25'h000_0001;
  assign p1_add_33413_comb = p1_umul_32948_comb[31:11] + p1_add_33354_comb;
  assign p1_add_33415_comb = p1_umul_33013_comb[31:1] + p1_umul_32986_comb[31:1];
  assign p1_add_33417_comb = p1_umul_32991_comb[31:7] + 25'h000_0001;
  assign p1_add_33419_comb = p1_umul_32952_comb[31:11] + p1_add_33360_comb;
  assign p1_add_33421_comb = p1_umul_33018_comb[31:1] + p1_umul_32992_comb[31:1];
  assign p1_add_33433_comb = p1_umul_33013_comb[31:7] + 25'h000_0001;
  assign p1_add_33435_comb = p1_umul_32986_comb[31:11] + p1_add_33354_comb;
  assign p1_add_33437_comb = p1_umul_32985_comb[31:3] + p1_umul_32948_comb[31:3];
  assign p1_add_33439_comb = p1_umul_33018_comb[31:7] + 25'h000_0001;
  assign p1_add_33441_comb = p1_umul_32992_comb[31:11] + p1_add_33360_comb;
  assign p1_add_33443_comb = p1_umul_32991_comb[31:3] + p1_umul_32952_comb[31:3];
  assign p1_add_33449_comb = p1_umul_33011_comb[31:7] + 25'h000_0001;
  assign p1_add_33451_comb = p1_add_33321_comb[26:6] + p1_add_33354_comb;
  assign p1_add_33453_comb = p1_umul_32985_comb[31:3] + p1_umul_32947_comb[31:3];
  assign p1_add_33455_comb = p1_umul_33016_comb[31:7] + 25'h000_0001;
  assign p1_add_33457_comb = p1_add_33322_comb[26:6] + p1_add_33360_comb;
  assign p1_add_33459_comb = p1_umul_32991_comb[31:3] + p1_umul_32951_comb[31:3];
  assign p1_add_33645_comb = p1_umul_33123_comb[31:7] + 25'h000_0001;
  assign p1_add_33647_comb = p1_umul_33076_comb[31:11] + p1_add_33610_comb;
  assign p1_add_33649_comb = p1_umul_33153_comb[31:1] + p1_umul_33124_comb[31:1];
  assign p1_add_33651_comb = p1_umul_33129_comb[31:7] + 25'h000_0001;
  assign p1_add_33653_comb = p1_umul_33080_comb[31:11] + p1_add_33616_comb;
  assign p1_add_33655_comb = p1_umul_33158_comb[31:1] + p1_umul_33130_comb[31:1];
  assign p1_add_33657_comb = p1_umul_33153_comb[31:7] + 25'h000_0001;
  assign p1_add_33659_comb = p1_umul_33124_comb[31:11] + p1_add_33610_comb;
  assign p1_add_33661_comb = p1_umul_33123_comb[31:3] + p1_umul_33076_comb[31:3];
  assign p1_add_33663_comb = p1_umul_33158_comb[31:7] + 25'h000_0001;
  assign p1_add_33665_comb = p1_umul_33130_comb[31:11] + p1_add_33616_comb;
  assign p1_add_33667_comb = p1_umul_33129_comb[31:3] + p1_umul_33080_comb[31:3];
  assign p1_add_33669_comb = p1_umul_33151_comb[31:7] + 25'h000_0001;
  assign p1_add_33671_comb = p1_add_33597_comb[26:6] + p1_add_33610_comb;
  assign p1_add_33673_comb = p1_umul_33123_comb[31:3] + p1_umul_33075_comb[31:3];
  assign p1_add_33675_comb = p1_umul_33156_comb[31:7] + 25'h000_0001;
  assign p1_add_33677_comb = p1_add_33598_comb[26:6] + p1_add_33616_comb;
  assign p1_add_33679_comb = p1_umul_33129_comb[31:3] + p1_umul_33079_comb[31:3];
  assign p1_add_32997_comb = p1_umul_32953_comb[31:3] + p1_umul_32954_comb[31:3];
  assign p1_add_32999_comb = p1_umul_32977_comb + p1_concat_32978_comb;
  assign p1_add_33000_comb = p1_umul_32979_comb + p1_umul_32920_comb;
  assign p1_add_33001_comb = p1_umul_32959_comb[31:3] + p1_umul_32960_comb[31:3];
  assign p1_add_33003_comb = p1_umul_32982_comb + p1_concat_32983_comb;
  assign p1_add_33004_comb = p1_umul_32984_comb + p1_umul_32924_comb;
  assign p1_add_33033_comb = p1_umul_32985_comb[31:3] + p1_umul_32986_comb[31:3];
  assign p1_add_33035_comb = p1_umul_33011_comb + p1_concat_33012_comb;
  assign p1_add_33036_comb = p1_umul_33013_comb + p1_umul_32948_comb;
  assign p1_add_33037_comb = p1_umul_32991_comb[31:3] + p1_umul_32992_comb[31:3];
  assign p1_add_33039_comb = p1_umul_33016_comb + p1_concat_33017_comb;
  assign p1_add_33040_comb = p1_umul_33018_comb + p1_umul_32952_comb;
  assign p1_add_33171_comb = p1_umul_33123_comb[31:3] + p1_umul_33124_comb[31:3];
  assign p1_add_33173_comb = p1_umul_33151_comb + p1_concat_33152_comb;
  assign p1_add_33174_comb = p1_umul_33153_comb + p1_umul_33076_comb;
  assign p1_add_33175_comb = p1_umul_33129_comb[31:3] + p1_umul_33130_comb[31:3];
  assign p1_add_33177_comb = p1_umul_33156_comb + p1_concat_33157_comb;
  assign p1_add_33178_comb = p1_umul_33158_comb + p1_umul_33080_comb;
  assign p1_sub_33345_comb = p1_umul_32953_comb - p1_umul_32977_comb;
  assign p1_sub_33348_comb = p1_umul_32959_comb - p1_umul_32982_comb;
  assign p1_concat_33366_comb = {p1_add_33221_comb, p1_umul_33168_comb[4:2]};
  assign p1_concat_33370_comb = {p1_add_33222_comb, p1_umul_33170_comb[4:2]};
  assign p1_sub_33473_comb = p1_umul_32985_comb - p1_umul_33011_comb;
  assign p1_sub_33476_comb = p1_umul_32991_comb - p1_umul_33016_comb;
  assign p1_concat_33486_comb = {p1_add_33321_comb, p1_umul_33218_comb[4:2]};
  assign p1_concat_33490_comb = {p1_add_33322_comb, p1_umul_33220_comb[4:2]};
  assign p1_sub_33683_comb = p1_umul_33123_comb - p1_umul_33151_comb;
  assign p1_sub_33686_comb = p1_umul_33129_comb - p1_umul_33156_comb;
  assign p1_concat_33692_comb = {p1_add_33597_comb, p1_umul_33520_comb[4:2]};
  assign p1_concat_33696_comb = {p1_add_33598_comb, p1_umul_33522_comb[4:2]};
  assign p1_add_33405_comb = p1_sub_33345_comb + p1_concat_32978_comb;
  assign p1_add_33406_comb = p1_add_33221_comb[26:2] + {p1_add_33248_comb, 4'h1};
  assign p1_add_33408_comb = p1_sub_33348_comb + p1_concat_32983_comb;
  assign p1_add_33409_comb = p1_add_33222_comb[26:2] + {p1_add_33254_comb, 4'h1};
  assign p1_add_33423_comb = {p1_add_33297_comb, p1_umul_32953_comb[6:3]} + {p1_add_33299_comb, p1_umul_32920_comb[10:3]};
  assign p1_add_33425_comb = p1_add_33301_comb[30:1] + p1_concat_33366_comb;
  assign p1_add_33428_comb = {p1_add_33303_comb, p1_umul_32959_comb[6:3]} + {p1_add_33305_comb, p1_umul_32924_comb[10:3]};
  assign p1_add_33430_comb = p1_add_33307_comb[30:1] + p1_concat_33370_comb;
  assign p1_add_33445_comb = {p1_add_33309_comb, p1_umul_32979_comb[6:1]} + {p1_add_33311_comb, p1_umul_32954_comb[10:1]};
  assign p1_add_33446_comb = {p1_add_33313_comb, p1_umul_32920_comb[2]} + p1_concat_33366_comb;
  assign p1_add_33447_comb = {p1_add_33315_comb, p1_umul_32984_comb[6:1]} + {p1_add_33317_comb, p1_umul_32960_comb[10:1]};
  assign p1_add_33448_comb = {p1_add_33319_comb, p1_umul_32924_comb[2]} + p1_concat_33370_comb;
  assign p1_add_33461_comb = {p1_add_33323_comb, p1_umul_32977_comb[6:2]} + {p1_add_33325_comb, p1_add_33221_comb[5:0], p1_umul_33168_comb[4:2]};
  assign p1_add_33463_comb = {p1_add_33327_comb, p1_umul_32919_comb[2]} + p1_umul_32920_comb[31:2];
  assign p1_add_33464_comb = {p1_add_33329_comb, p1_umul_32982_comb[6:2]} + {p1_add_33331_comb, p1_add_33222_comb[5:0], p1_umul_33170_comb[4:2]};
  assign p1_add_33466_comb = {p1_add_33333_comb, p1_umul_32923_comb[2]} + p1_umul_32924_comb[31:2];
  assign p1_add_33523_comb = p1_sub_33473_comb + p1_concat_33012_comb;
  assign p1_add_33524_comb = p1_add_33321_comb[26:2] + {p1_add_33354_comb, 4'h1};
  assign p1_add_33526_comb = p1_sub_33476_comb + p1_concat_33017_comb;
  assign p1_add_33527_comb = p1_add_33322_comb[26:2] + {p1_add_33360_comb, 4'h1};
  assign p1_add_33531_comb = {p1_add_33411_comb, p1_umul_32985_comb[6:3]} + {p1_add_33413_comb, p1_umul_32948_comb[10:3]};
  assign p1_add_33533_comb = p1_add_33415_comb[30:1] + p1_concat_33486_comb;
  assign p1_add_33536_comb = {p1_add_33417_comb, p1_umul_32991_comb[6:3]} + {p1_add_33419_comb, p1_umul_32952_comb[10:3]};
  assign p1_add_33538_comb = p1_add_33421_comb[30:1] + p1_concat_33490_comb;
  assign p1_add_33543_comb = {p1_add_33433_comb, p1_umul_33013_comb[6:1]} + {p1_add_33435_comb, p1_umul_32986_comb[10:1]};
  assign p1_add_33544_comb = {p1_add_33437_comb, p1_umul_32948_comb[2]} + p1_concat_33486_comb;
  assign p1_add_33545_comb = {p1_add_33439_comb, p1_umul_33018_comb[6:1]} + {p1_add_33441_comb, p1_umul_32992_comb[10:1]};
  assign p1_add_33546_comb = {p1_add_33443_comb, p1_umul_32952_comb[2]} + p1_concat_33490_comb;
  assign p1_add_33549_comb = {p1_add_33449_comb, p1_umul_33011_comb[6:2]} + {p1_add_33451_comb, p1_add_33321_comb[5:0], p1_umul_33218_comb[4:2]};
  assign p1_add_33551_comb = {p1_add_33453_comb, p1_umul_32947_comb[2]} + p1_umul_32948_comb[31:2];
  assign p1_add_33552_comb = {p1_add_33455_comb, p1_umul_33016_comb[6:2]} + {p1_add_33457_comb, p1_add_33322_comb[5:0], p1_umul_33220_comb[4:2]};
  assign p1_add_33554_comb = {p1_add_33459_comb, p1_umul_32951_comb[2]} + p1_umul_32952_comb[31:2];
  assign p1_add_33713_comb = p1_sub_33683_comb + p1_concat_33152_comb;
  assign p1_add_33714_comb = p1_add_33597_comb[26:2] + {p1_add_33610_comb, 4'h1};
  assign p1_add_33716_comb = p1_sub_33686_comb + p1_concat_33157_comb;
  assign p1_add_33717_comb = p1_add_33598_comb[26:2] + {p1_add_33616_comb, 4'h1};
  assign p1_add_33719_comb = {p1_add_33645_comb, p1_umul_33123_comb[6:3]} + {p1_add_33647_comb, p1_umul_33076_comb[10:3]};
  assign p1_add_33721_comb = p1_add_33649_comb[30:1] + p1_concat_33692_comb;
  assign p1_add_33724_comb = {p1_add_33651_comb, p1_umul_33129_comb[6:3]} + {p1_add_33653_comb, p1_umul_33080_comb[10:3]};
  assign p1_add_33726_comb = p1_add_33655_comb[30:1] + p1_concat_33696_comb;
  assign p1_add_33729_comb = {p1_add_33657_comb, p1_umul_33153_comb[6:1]} + {p1_add_33659_comb, p1_umul_33124_comb[10:1]};
  assign p1_add_33730_comb = {p1_add_33661_comb, p1_umul_33076_comb[2]} + p1_concat_33692_comb;
  assign p1_add_33731_comb = {p1_add_33663_comb, p1_umul_33158_comb[6:1]} + {p1_add_33665_comb, p1_umul_33130_comb[10:1]};
  assign p1_add_33732_comb = {p1_add_33667_comb, p1_umul_33080_comb[2]} + p1_concat_33696_comb;
  assign p1_add_33733_comb = {p1_add_33669_comb, p1_umul_33151_comb[6:2]} + {p1_add_33671_comb, p1_add_33597_comb[5:0], p1_umul_33520_comb[4:2]};
  assign p1_add_33735_comb = {p1_add_33673_comb, p1_umul_33075_comb[2]} + p1_umul_33076_comb[31:2];
  assign p1_add_33736_comb = {p1_add_33675_comb, p1_umul_33156_comb[6:2]} + {p1_add_33677_comb, p1_add_33598_comb[5:0], p1_umul_33522_comb[4:2]};
  assign p1_add_33738_comb = {p1_add_33679_comb, p1_umul_33079_comb[2]} + p1_umul_33080_comb[31:2];
  assign p1_add_33029_comb = p1_add_32997_comb + p1_umul_32953_comb[31:3];
  assign p1_add_33031_comb = p1_add_33001_comb + p1_umul_32959_comb[31:3];
  assign p1_add_33041_comb = {p1_add_32997_comb, p1_umul_32954_comb[2:1]} + p1_add_32999_comb[31:1];
  assign p1_add_33043_comb = p1_add_33000_comb[31:3] + p1_umul_32953_comb[31:3];
  assign p1_add_33045_comb = {p1_add_33001_comb, p1_umul_32960_comb[2:1]} + p1_add_33003_comb[31:1];
  assign p1_add_33047_comb = p1_add_33004_comb[31:3] + p1_umul_32959_comb[31:3];
  assign p1_add_33081_comb = p1_add_33033_comb + p1_umul_32985_comb[31:3];
  assign p1_add_33083_comb = p1_add_33037_comb + p1_umul_32991_comb[31:3];
  assign p1_add_33087_comb = {p1_add_33033_comb, p1_umul_32986_comb[2:1]} + p1_add_33035_comb[31:1];
  assign p1_add_33089_comb = p1_add_33036_comb[31:3] + p1_umul_32985_comb[31:3];
  assign p1_add_33091_comb = {p1_add_33037_comb, p1_umul_32992_comb[2:1]} + p1_add_33039_comb[31:1];
  assign p1_add_33093_comb = p1_add_33040_comb[31:3] + p1_umul_32991_comb[31:3];
  assign p1_add_33223_comb = p1_add_33171_comb + p1_umul_33123_comb[31:3];
  assign p1_add_33225_comb = p1_add_33175_comb + p1_umul_33129_comb[31:3];
  assign p1_add_33227_comb = {p1_add_33171_comb, p1_umul_33124_comb[2:1]} + p1_add_33173_comb[31:1];
  assign p1_add_33229_comb = p1_add_33174_comb[31:3] + p1_umul_33123_comb[31:3];
  assign p1_add_33231_comb = {p1_add_33175_comb, p1_umul_33130_comb[2:1]} + p1_add_33177_comb[31:1];
  assign p1_add_33233_comb = p1_add_33178_comb[31:3] + p1_umul_33129_comb[31:3];
  assign p1_add_33059_comb = p1_add_32999_comb + p1_add_33000_comb;
  assign p1_add_33061_comb = p1_add_33003_comb + p1_add_33004_comb;
  assign p1_add_33111_comb = p1_add_33035_comb + p1_add_33036_comb;
  assign p1_add_33113_comb = p1_add_33039_comb + p1_add_33040_comb;
  assign p1_add_33277_comb = p1_add_33173_comb + p1_add_33174_comb;
  assign p1_add_33279_comb = p1_add_33177_comb + p1_add_33178_comb;
  assign p1_add_33529_comb = p1_add_33405_comb[31:2] + {p1_add_33406_comb, p1_add_33221_comb[1:0], p1_umul_33168_comb[4:2]};
  assign p1_add_33530_comb = p1_add_33408_comb[31:2] + {p1_add_33409_comb, p1_add_33222_comb[1:0], p1_umul_33170_comb[4:2]};
  assign p1_sub_33541_comb = {p1_add_33423_comb, p1_umul_32920_comb[2:0]} - {p1_add_33425_comb, p1_add_33301_comb[0], p1_umul_32979_comb[0]};
  assign p1_sub_33542_comb = {p1_add_33428_comb, p1_umul_32924_comb[2:0]} - {p1_add_33430_comb, p1_add_33307_comb[0], p1_umul_32984_comb[0]};
  assign p1_sub_33547_comb = {p1_add_33445_comb, p1_umul_32979_comb[0]} - {p1_add_33446_comb, p1_umul_32920_comb[1:0]};
  assign p1_sub_33548_comb = {p1_add_33447_comb, p1_umul_32984_comb[0]} - {p1_add_33448_comb, p1_umul_32924_comb[1:0]};
  assign p1_sub_33555_comb = {p1_add_33461_comb, p1_umul_32977_comb[1:0]} - {p1_add_33463_comb, p1_umul_32920_comb[1:0]};
  assign p1_sub_33556_comb = {p1_add_33464_comb, p1_umul_32982_comb[1:0]} - {p1_add_33466_comb, p1_umul_32924_comb[1:0]};
  assign p1_add_33599_comb = p1_add_33523_comb[31:2] + {p1_add_33524_comb, p1_add_33321_comb[1:0], p1_umul_33218_comb[4:2]};
  assign p1_add_33600_comb = p1_add_33526_comb[31:2] + {p1_add_33527_comb, p1_add_33322_comb[1:0], p1_umul_33220_comb[4:2]};
  assign p1_sub_33601_comb = {p1_add_33531_comb, p1_umul_32948_comb[2:0]} - {p1_add_33533_comb, p1_add_33415_comb[0], p1_umul_33013_comb[0]};
  assign p1_sub_33602_comb = {p1_add_33536_comb, p1_umul_32952_comb[2:0]} - {p1_add_33538_comb, p1_add_33421_comb[0], p1_umul_33018_comb[0]};
  assign p1_sub_33603_comb = {p1_add_33543_comb, p1_umul_33013_comb[0]} - {p1_add_33544_comb, p1_umul_32948_comb[1:0]};
  assign p1_sub_33604_comb = {p1_add_33545_comb, p1_umul_33018_comb[0]} - {p1_add_33546_comb, p1_umul_32952_comb[1:0]};
  assign p1_sub_33605_comb = {p1_add_33549_comb, p1_umul_33011_comb[1:0]} - {p1_add_33551_comb, p1_umul_32948_comb[1:0]};
  assign p1_sub_33606_comb = {p1_add_33552_comb, p1_umul_33016_comb[1:0]} - {p1_add_33554_comb, p1_umul_32952_comb[1:0]};
  assign p1_add_33759_comb = p1_add_33713_comb[31:2] + {p1_add_33714_comb, p1_add_33597_comb[1:0], p1_umul_33520_comb[4:2]};
  assign p1_add_33760_comb = p1_add_33716_comb[31:2] + {p1_add_33717_comb, p1_add_33598_comb[1:0], p1_umul_33522_comb[4:2]};
  assign p1_sub_33761_comb = {p1_add_33719_comb, p1_umul_33076_comb[2:0]} - {p1_add_33721_comb, p1_add_33649_comb[0], p1_umul_33153_comb[0]};
  assign p1_sub_33762_comb = {p1_add_33724_comb, p1_umul_33080_comb[2:0]} - {p1_add_33726_comb, p1_add_33655_comb[0], p1_umul_33158_comb[0]};
  assign p1_sub_33763_comb = {p1_add_33729_comb, p1_umul_33153_comb[0]} - {p1_add_33730_comb, p1_umul_33076_comb[1:0]};
  assign p1_sub_33764_comb = {p1_add_33731_comb, p1_umul_33158_comb[0]} - {p1_add_33732_comb, p1_umul_33080_comb[1:0]};
  assign p1_sub_33765_comb = {p1_add_33733_comb, p1_umul_33151_comb[1:0]} - {p1_add_33735_comb, p1_umul_33076_comb[1:0]};
  assign p1_sub_33766_comb = {p1_add_33736_comb, p1_umul_33156_comb[1:0]} - {p1_add_33738_comb, p1_umul_33080_comb[1:0]};
  assign p1_sub_33085_comb = p1_add_33059_comb - {p1_add_33029_comb, p1_umul_32954_comb[2:0]};
  assign p1_sub_33086_comb = p1_add_33061_comb - {p1_add_33031_comb, p1_umul_32960_comb[2:0]};
  assign p1_sub_33095_comb = {p1_add_33041_comb, p1_add_32999_comb[0]} - {p1_add_33043_comb, p1_add_33000_comb[2:0]};
  assign p1_sub_33096_comb = {p1_add_33045_comb, p1_add_33003_comb[0]} - {p1_add_33047_comb, p1_add_33004_comb[2:0]};
  assign p1_sub_33135_comb = p1_add_33111_comb - {p1_add_33081_comb, p1_umul_32986_comb[2:0]};
  assign p1_sub_33136_comb = p1_add_33113_comb - {p1_add_33083_comb, p1_umul_32992_comb[2:0]};
  assign p1_sub_33137_comb = {p1_add_33087_comb, p1_add_33035_comb[0]} - {p1_add_33089_comb, p1_add_33036_comb[2:0]};
  assign p1_sub_33138_comb = {p1_add_33091_comb, p1_add_33039_comb[0]} - {p1_add_33093_comb, p1_add_33040_comb[2:0]};
  assign p1_array_index_33203_comb = p0_f[6'h01];
  assign p1_array_index_33204_comb = p0_f[6'h07];
  assign p1_array_index_33237_comb = p0_f[6'h21];
  assign p1_array_index_33238_comb = p0_f[6'h27];
  assign p1_array_index_33285_comb = p0_f[6'h05];
  assign p1_array_index_33286_comb = p0_f[6'h03];
  assign p1_sub_33335_comb = p1_add_33277_comb - {p1_add_33223_comb, p1_umul_33124_comb[2:0]};
  assign p1_sub_33336_comb = p1_add_33279_comb - {p1_add_33225_comb, p1_umul_33130_comb[2:0]};
  assign p1_sub_33337_comb = {p1_add_33227_comb, p1_add_33173_comb[0]} - {p1_add_33229_comb, p1_add_33174_comb[2:0]};
  assign p1_sub_33338_comb = {p1_add_33231_comb, p1_add_33177_comb[0]} - {p1_add_33233_comb, p1_add_33178_comb[2:0]};
  assign p1_array_index_33343_comb = p0_f[6'h25];
  assign p1_array_index_33344_comb = p0_f[6'h23];
  assign p1_bit_slice_33571_comb = p1_add_33529_comb[29:6];
  assign p1_bit_slice_33572_comb = p1_add_33530_comb[29:6];
  assign p1_bit_slice_33577_comb = p1_sub_33541_comb[31:8];
  assign p1_bit_slice_33578_comb = p1_sub_33542_comb[31:8];
  assign p1_bit_slice_33583_comb = p1_sub_33547_comb[31:8];
  assign p1_bit_slice_33584_comb = p1_sub_33548_comb[31:8];
  assign p1_bit_slice_33589_comb = p1_sub_33555_comb[31:8];
  assign p1_bit_slice_33590_comb = p1_sub_33556_comb[31:8];
  assign p1_bit_slice_33635_comb = p1_add_33599_comb[29:6];
  assign p1_bit_slice_33636_comb = p1_add_33600_comb[29:6];
  assign p1_bit_slice_33637_comb = p1_sub_33601_comb[31:8];
  assign p1_bit_slice_33638_comb = p1_sub_33602_comb[31:8];
  assign p1_bit_slice_33639_comb = p1_sub_33603_comb[31:8];
  assign p1_bit_slice_33640_comb = p1_sub_33604_comb[31:8];
  assign p1_bit_slice_33641_comb = p1_sub_33605_comb[31:8];
  assign p1_bit_slice_33642_comb = p1_sub_33606_comb[31:8];
  assign p1_array_index_33709_comb = p0_f[6'h02];
  assign p1_array_index_33710_comb = p0_f[6'h06];
  assign p1_array_index_33739_comb = p0_f[6'h22];
  assign p1_array_index_33740_comb = p0_f[6'h26];
  assign p1_bit_slice_33771_comb = p1_add_33759_comb[29:6];
  assign p1_bit_slice_33772_comb = p1_add_33760_comb[29:6];
  assign p1_bit_slice_33773_comb = p1_sub_33761_comb[31:8];
  assign p1_bit_slice_33774_comb = p1_sub_33762_comb[31:8];
  assign p1_bit_slice_33775_comb = p1_sub_33763_comb[31:8];
  assign p1_bit_slice_33776_comb = p1_sub_33764_comb[31:8];
  assign p1_bit_slice_33777_comb = p1_sub_33765_comb[31:8];
  assign p1_bit_slice_33778_comb = p1_sub_33766_comb[31:8];
  assign p1_bit_slice_33779_comb = p0_f[6'h04][20:0];
  assign p1_bit_slice_33780_comb = p0_f[6'h00][20:0];
  assign p1_bit_slice_33783_comb = p0_f[6'h24][20:0];
  assign p1_bit_slice_33784_comb = p0_f[6'h20][20:0];
  assign p1_umul_33207_comb = umul32b_32b_x_12b(p1_array_index_33120_comb, 12'hec8);
  assign p1_umul_33208_comb = umul32b_32b_x_12b(p1_array_index_33122_comb, 12'hec8);
  assign p1_umul_33291_comb = umul32b_32b_x_12b(p1_array_index_33164_comb, 12'hec8);
  assign p1_umul_33292_comb = umul32b_32b_x_12b(p1_array_index_33166_comb, 12'hec8);
  assign p1_umul_33591_comb = umul32b_32b_x_12b(p1_array_index_33400_comb, 12'hec8);
  assign p1_umul_33592_comb = umul32b_32b_x_12b(p1_array_index_33402_comb, 12'hec8);

  // Registers for pipe stage 1:
  reg [31:0] p1_sub_33085;
  reg [31:0] p1_sub_33086;
  reg [31:0] p1_sub_33095;
  reg [31:0] p1_sub_33096;
  reg [31:0] p1_sub_33135;
  reg [31:0] p1_sub_33136;
  reg [31:0] p1_sub_33137;
  reg [31:0] p1_sub_33138;
  reg [31:0] p1_array_index_33203;
  reg [31:0] p1_array_index_33204;
  reg [20:0] p1_bit_slice_33213;
  reg [20:0] p1_bit_slice_33214;
  reg [20:0] p1_bit_slice_33215;
  reg [20:0] p1_bit_slice_33216;
  reg [31:0] p1_array_index_33237;
  reg [31:0] p1_array_index_33238;
  reg [31:0] p1_array_index_33285;
  reg [31:0] p1_array_index_33286;
  reg [20:0] p1_bit_slice_33293;
  reg [20:0] p1_bit_slice_33294;
  reg [20:0] p1_bit_slice_33295;
  reg [20:0] p1_bit_slice_33296;
  reg [31:0] p1_sub_33335;
  reg [31:0] p1_sub_33336;
  reg [31:0] p1_sub_33337;
  reg [31:0] p1_sub_33338;
  reg [31:0] p1_array_index_33343;
  reg [31:0] p1_array_index_33344;
  reg [23:0] p1_bit_slice_33571;
  reg [23:0] p1_bit_slice_33572;
  reg [23:0] p1_bit_slice_33577;
  reg [23:0] p1_bit_slice_33578;
  reg [23:0] p1_bit_slice_33583;
  reg [23:0] p1_bit_slice_33584;
  reg [23:0] p1_bit_slice_33589;
  reg [23:0] p1_bit_slice_33590;
  reg [20:0] p1_bit_slice_33593;
  reg [20:0] p1_bit_slice_33594;
  reg [20:0] p1_bit_slice_33595;
  reg [20:0] p1_bit_slice_33596;
  reg [23:0] p1_bit_slice_33635;
  reg [23:0] p1_bit_slice_33636;
  reg [23:0] p1_bit_slice_33637;
  reg [23:0] p1_bit_slice_33638;
  reg [23:0] p1_bit_slice_33639;
  reg [23:0] p1_bit_slice_33640;
  reg [23:0] p1_bit_slice_33641;
  reg [23:0] p1_bit_slice_33642;
  reg [31:0] p1_array_index_33709;
  reg [31:0] p1_array_index_33710;
  reg [31:0] p1_array_index_33739;
  reg [31:0] p1_array_index_33740;
  reg [23:0] p1_bit_slice_33771;
  reg [23:0] p1_bit_slice_33772;
  reg [23:0] p1_bit_slice_33773;
  reg [23:0] p1_bit_slice_33774;
  reg [23:0] p1_bit_slice_33775;
  reg [23:0] p1_bit_slice_33776;
  reg [23:0] p1_bit_slice_33777;
  reg [23:0] p1_bit_slice_33778;
  reg [20:0] p1_bit_slice_33779;
  reg [20:0] p1_bit_slice_33780;
  reg [20:0] p1_bit_slice_33783;
  reg [20:0] p1_bit_slice_33784;
  reg [31:0] p1_umul_33168;
  reg [31:0] p1_umul_33170;
  reg [31:0] p1_umul_33207;
  reg [31:0] p1_umul_33208;
  reg [31:0] p1_umul_33218;
  reg [31:0] p1_umul_33220;
  reg [31:0] p1_umul_33291;
  reg [31:0] p1_umul_33292;
  reg [31:0] p1_umul_33520;
  reg [31:0] p1_umul_33522;
  reg [31:0] p1_umul_33591;
  reg [31:0] p1_umul_33592;
  always_ff @ (posedge clk) begin
    p1_sub_33085 <= p1_sub_33085_comb;
    p1_sub_33086 <= p1_sub_33086_comb;
    p1_sub_33095 <= p1_sub_33095_comb;
    p1_sub_33096 <= p1_sub_33096_comb;
    p1_sub_33135 <= p1_sub_33135_comb;
    p1_sub_33136 <= p1_sub_33136_comb;
    p1_sub_33137 <= p1_sub_33137_comb;
    p1_sub_33138 <= p1_sub_33138_comb;
    p1_array_index_33203 <= p1_array_index_33203_comb;
    p1_array_index_33204 <= p1_array_index_33204_comb;
    p1_bit_slice_33213 <= p1_bit_slice_33213_comb;
    p1_bit_slice_33214 <= p1_bit_slice_33214_comb;
    p1_bit_slice_33215 <= p1_bit_slice_33215_comb;
    p1_bit_slice_33216 <= p1_bit_slice_33216_comb;
    p1_array_index_33237 <= p1_array_index_33237_comb;
    p1_array_index_33238 <= p1_array_index_33238_comb;
    p1_array_index_33285 <= p1_array_index_33285_comb;
    p1_array_index_33286 <= p1_array_index_33286_comb;
    p1_bit_slice_33293 <= p1_bit_slice_33293_comb;
    p1_bit_slice_33294 <= p1_bit_slice_33294_comb;
    p1_bit_slice_33295 <= p1_bit_slice_33295_comb;
    p1_bit_slice_33296 <= p1_bit_slice_33296_comb;
    p1_sub_33335 <= p1_sub_33335_comb;
    p1_sub_33336 <= p1_sub_33336_comb;
    p1_sub_33337 <= p1_sub_33337_comb;
    p1_sub_33338 <= p1_sub_33338_comb;
    p1_array_index_33343 <= p1_array_index_33343_comb;
    p1_array_index_33344 <= p1_array_index_33344_comb;
    p1_bit_slice_33571 <= p1_bit_slice_33571_comb;
    p1_bit_slice_33572 <= p1_bit_slice_33572_comb;
    p1_bit_slice_33577 <= p1_bit_slice_33577_comb;
    p1_bit_slice_33578 <= p1_bit_slice_33578_comb;
    p1_bit_slice_33583 <= p1_bit_slice_33583_comb;
    p1_bit_slice_33584 <= p1_bit_slice_33584_comb;
    p1_bit_slice_33589 <= p1_bit_slice_33589_comb;
    p1_bit_slice_33590 <= p1_bit_slice_33590_comb;
    p1_bit_slice_33593 <= p1_bit_slice_33593_comb;
    p1_bit_slice_33594 <= p1_bit_slice_33594_comb;
    p1_bit_slice_33595 <= p1_bit_slice_33595_comb;
    p1_bit_slice_33596 <= p1_bit_slice_33596_comb;
    p1_bit_slice_33635 <= p1_bit_slice_33635_comb;
    p1_bit_slice_33636 <= p1_bit_slice_33636_comb;
    p1_bit_slice_33637 <= p1_bit_slice_33637_comb;
    p1_bit_slice_33638 <= p1_bit_slice_33638_comb;
    p1_bit_slice_33639 <= p1_bit_slice_33639_comb;
    p1_bit_slice_33640 <= p1_bit_slice_33640_comb;
    p1_bit_slice_33641 <= p1_bit_slice_33641_comb;
    p1_bit_slice_33642 <= p1_bit_slice_33642_comb;
    p1_array_index_33709 <= p1_array_index_33709_comb;
    p1_array_index_33710 <= p1_array_index_33710_comb;
    p1_array_index_33739 <= p1_array_index_33739_comb;
    p1_array_index_33740 <= p1_array_index_33740_comb;
    p1_bit_slice_33771 <= p1_bit_slice_33771_comb;
    p1_bit_slice_33772 <= p1_bit_slice_33772_comb;
    p1_bit_slice_33773 <= p1_bit_slice_33773_comb;
    p1_bit_slice_33774 <= p1_bit_slice_33774_comb;
    p1_bit_slice_33775 <= p1_bit_slice_33775_comb;
    p1_bit_slice_33776 <= p1_bit_slice_33776_comb;
    p1_bit_slice_33777 <= p1_bit_slice_33777_comb;
    p1_bit_slice_33778 <= p1_bit_slice_33778_comb;
    p1_bit_slice_33779 <= p1_bit_slice_33779_comb;
    p1_bit_slice_33780 <= p1_bit_slice_33780_comb;
    p1_bit_slice_33783 <= p1_bit_slice_33783_comb;
    p1_bit_slice_33784 <= p1_bit_slice_33784_comb;
    p1_umul_33168 <= p1_umul_33168_comb;
    p1_umul_33170 <= p1_umul_33170_comb;
    p1_umul_33207 <= p1_umul_33207_comb;
    p1_umul_33208 <= p1_umul_33208_comb;
    p1_umul_33218 <= p1_umul_33218_comb;
    p1_umul_33220 <= p1_umul_33220_comb;
    p1_umul_33291 <= p1_umul_33291_comb;
    p1_umul_33292 <= p1_umul_33292_comb;
    p1_umul_33520 <= p1_umul_33520_comb;
    p1_umul_33522 <= p1_umul_33522_comb;
    p1_umul_33591 <= p1_umul_33591_comb;
    p1_umul_33592 <= p1_umul_33592_comb;
  end

  // ===== Pipe stage 2:
  wire [31:0] p2_umul_33941_comb;
  wire [31:0] p2_umul_33942_comb;
  wire [31:0] p2_umul_33943_comb;
  wire [31:0] p2_umul_33944_comb;
  wire [31:0] p2_umul_33957_comb;
  wire [31:0] p2_umul_33958_comb;
  wire [24:0] p2_add_33959_comb;
  wire [24:0] p2_add_33960_comb;
  wire [31:0] p2_umul_33961_comb;
  wire [31:0] p2_umul_33962_comb;
  wire [24:0] p2_add_33963_comb;
  wire [24:0] p2_add_33964_comb;
  wire [31:0] p2_add_34598_comb;
  wire [23:0] p2_bit_slice_33969_comb;
  wire [23:0] p2_bit_slice_33970_comb;
  wire [23:0] p2_bit_slice_33975_comb;
  wire [23:0] p2_bit_slice_33976_comb;
  wire [31:0] p2_umul_34686_comb;
  wire [31:0] p2_umul_34687_comb;
  wire [31:0] p2_add_34689_comb;
  wire [24:0] p2_add_33977_comb;
  wire [24:0] p2_add_33978_comb;
  wire [31:0] p2_sign_ext_33979_comb;
  wire [31:0] p2_sign_ext_33980_comb;
  wire [24:0] p2_add_33981_comb;
  wire [24:0] p2_add_33982_comb;
  wire [31:0] p2_sign_ext_33983_comb;
  wire [31:0] p2_sign_ext_33984_comb;
  wire [31:0] p2_add_34057_comb;
  wire [31:0] p2_add_33986_comb;
  wire [31:0] p2_umul_34752_comb;
  wire [31:0] p2_umul_34753_comb;
  wire [23:0] p2_bit_slice_33988_comb;
  wire [23:0] p2_bit_slice_33989_comb;
  wire [23:0] p2_bit_slice_33996_comb;
  wire [23:0] p2_bit_slice_33997_comb;
  wire [31:0] p2_umul_34112_comb;
  wire [31:0] p2_umul_34021_comb;
  wire [31:0] p2_umul_34199_comb;
  wire [31:0] p2_umul_34113_comb;
  wire [31:0] p2_umul_34197_comb;
  wire [26:0] p2_add_34796_comb;
  wire [31:0] p2_umul_34020_comb;
  wire [31:0] p2_add_34118_comb;
  wire [31:0] p2_add_34023_comb;
  wire [31:0] p2_sign_ext_34025_comb;
  wire [31:0] p2_sign_ext_34026_comb;
  wire [24:0] p2_add_34027_comb;
  wire [20:0] p2_add_34029_comb;
  wire [24:0] p2_add_34031_comb;
  wire [20:0] p2_add_34033_comb;
  wire [31:0] p2_sign_ext_34035_comb;
  wire [31:0] p2_sign_ext_34036_comb;
  wire [24:0] p2_add_34037_comb;
  wire [20:0] p2_add_34039_comb;
  wire [24:0] p2_add_34041_comb;
  wire [20:0] p2_add_34043_comb;
  wire [24:0] p2_add_34045_comb;
  wire [29:0] p2_add_34046_comb;
  wire [24:0] p2_add_34047_comb;
  wire [29:0] p2_add_34048_comb;
  wire [24:0] p2_add_34049_comb;
  wire [28:0] p2_add_34050_comb;
  wire [24:0] p2_add_34051_comb;
  wire [28:0] p2_add_34052_comb;
  wire [31:0] p2_sign_ext_34831_comb;
  wire [31:0] p2_sign_ext_34832_comb;
  wire [20:0] p2_add_34841_comb;
  wire [31:0] p2_sign_ext_34833_comb;
  wire [31:0] p2_sign_ext_34834_comb;
  wire [31:0] p2_sign_ext_34835_comb;
  wire [31:0] p2_sign_ext_34836_comb;
  wire [31:0] p2_umul_34200_comb;
  wire [31:0] p2_umul_34063_comb;
  wire [31:0] p2_umul_34250_comb;
  wire [31:0] p2_umul_34201_comb;
  wire [31:0] p2_umul_34248_comb;
  wire [26:0] p2_add_34852_comb;
  wire [31:0] p2_umul_34062_comb;
  wire [31:0] p2_sign_ext_34347_comb;
  wire [31:0] p2_sign_ext_34348_comb;
  wire [31:0] p2_sign_ext_34357_comb;
  wire [31:0] p2_sign_ext_34358_comb;
  wire [31:0] p2_sign_ext_34359_comb;
  wire [31:0] p2_sign_ext_34360_comb;
  wire [31:0] p2_sign_ext_34369_comb;
  wire [31:0] p2_sign_ext_34370_comb;
  wire [31:0] p2_add_34869_comb;
  wire [24:0] p2_add_34876_comb;
  wire [20:0] p2_add_34878_comb;
  wire [30:0] p2_add_34880_comb;
  wire [31:0] p2_add_34871_comb;
  wire [24:0] p2_add_34888_comb;
  wire [20:0] p2_add_34890_comb;
  wire [28:0] p2_add_34892_comb;
  wire [31:0] p2_add_34873_comb;
  wire [24:0] p2_add_34898_comb;
  wire [20:0] p2_add_34900_comb;
  wire [28:0] p2_add_34902_comb;
  wire [20:0] p2_add_34885_comb;
  wire [31:0] p2_add_34409_comb;
  wire [31:0] p2_add_34419_comb;
  wire [31:0] p2_add_34421_comb;
  wire [31:0] p2_add_34431_comb;
  wire [24:0] p2_add_34123_comb;
  wire [20:0] p2_add_34125_comb;
  wire [24:0] p2_add_34127_comb;
  wire [20:0] p2_add_34129_comb;
  wire [29:0] p2_add_34131_comb;
  wire [20:0] p2_add_34133_comb;
  wire [29:0] p2_add_34135_comb;
  wire [20:0] p2_add_34137_comb;
  wire [24:0] p2_add_34139_comb;
  wire [20:0] p2_add_34141_comb;
  wire [24:0] p2_add_34143_comb;
  wire [20:0] p2_add_34145_comb;
  wire [28:0] p2_add_34147_comb;
  wire [20:0] p2_add_34149_comb;
  wire [28:0] p2_add_34151_comb;
  wire [20:0] p2_add_34153_comb;
  wire [24:0] p2_add_34155_comb;
  wire [29:0] p2_add_34156_comb;
  wire [24:0] p2_add_34157_comb;
  wire [29:0] p2_add_34158_comb;
  wire [20:0] p2_add_34159_comb;
  wire [20:0] p2_add_34162_comb;
  wire [20:0] p2_add_34165_comb;
  wire [20:0] p2_add_34168_comb;
  wire [24:0] p2_add_34171_comb;
  wire [28:0] p2_add_34172_comb;
  wire [24:0] p2_add_34173_comb;
  wire [28:0] p2_add_34174_comb;
  wire [20:0] p2_add_34175_comb;
  wire [20:0] p2_add_34178_comb;
  wire [20:0] p2_add_34181_comb;
  wire [20:0] p2_add_34184_comb;
  wire [31:0] p2_umul_34108_comb;
  wire [31:0] p2_umul_34109_comb;
  wire [31:0] p2_umul_34110_comb;
  wire [31:0] p2_umul_34111_comb;
  wire [31:0] p2_umul_34916_comb;
  wire [29:0] p2_concat_34926_comb;
  wire [31:0] p2_umul_34917_comb;
  wire [31:0] p2_umul_34918_comb;
  wire [24:0] p2_add_34927_comb;
  wire [20:0] p2_add_34929_comb;
  wire [30:0] p2_add_34931_comb;
  wire [24:0] p2_add_34936_comb;
  wire [20:0] p2_add_34938_comb;
  wire [28:0] p2_add_34940_comb;
  wire [24:0] p2_add_34945_comb;
  wire [20:0] p2_add_34947_comb;
  wire [28:0] p2_add_34949_comb;
  wire [31:0] p2_sign_ext_34465_comb;
  wire [31:0] p2_sign_ext_34466_comb;
  wire [31:0] p2_umul_34467_comb;
  wire [31:0] p2_sign_ext_34474_comb;
  wire [31:0] p2_sign_ext_34475_comb;
  wire [31:0] p2_umul_34476_comb;
  wire [31:0] p2_sign_ext_34477_comb;
  wire [31:0] p2_sign_ext_34478_comb;
  wire [31:0] p2_umul_34479_comb;
  wire [31:0] p2_sign_ext_34486_comb;
  wire [31:0] p2_sign_ext_34487_comb;
  wire [31:0] p2_umul_34488_comb;
  wire [28:0] p2_add_34971_comb;
  wire [29:0] p2_add_34973_comb;
  wire [30:0] p2_add_34980_comb;
  wire [29:0] p2_add_34981_comb;
  wire [29:0] p2_add_34985_comb;
  wire [29:0] p2_add_34987_comb;
  wire [29:0] p2_concat_34979_comb;
  wire [31:0] p2_add_34512_comb;
  wire [31:0] p2_add_34527_comb;
  wire [31:0] p2_add_34532_comb;
  wire [31:0] p2_add_34547_comb;
  wire [29:0] p2_add_34251_comb;
  wire [20:0] p2_add_34253_comb;
  wire [29:0] p2_add_34255_comb;
  wire [20:0] p2_add_34257_comb;
  wire [31:0] p2_sub_34259_comb;
  wire [31:0] p2_sub_34260_comb;
  wire [28:0] p2_add_34261_comb;
  wire [20:0] p2_add_34263_comb;
  wire [28:0] p2_add_34265_comb;
  wire [20:0] p2_add_34267_comb;
  wire [31:0] p2_sub_34269_comb;
  wire [31:0] p2_sub_34270_comb;
  wire [20:0] p2_add_34271_comb;
  wire [20:0] p2_add_34274_comb;
  wire [20:0] p2_add_34277_comb;
  wire [20:0] p2_add_34280_comb;
  wire [31:0] p2_sub_34283_comb;
  wire [31:0] p2_sub_34284_comb;
  wire [20:0] p2_add_34285_comb;
  wire [20:0] p2_add_34288_comb;
  wire [20:0] p2_add_34291_comb;
  wire [20:0] p2_add_34294_comb;
  wire [31:0] p2_sub_34297_comb;
  wire [31:0] p2_sub_34298_comb;
  wire [24:0] p2_add_34238_comb;
  wire [24:0] p2_add_34239_comb;
  wire [24:0] p2_add_34240_comb;
  wire [24:0] p2_add_34241_comb;
  wire [31:0] p2_umul_35058_comb;
  wire [29:0] p2_add_34997_comb;
  wire [31:0] p2_umul_35059_comb;
  wire [29:0] p2_add_35002_comb;
  wire [31:0] p2_umul_35060_comb;
  wire [29:0] p2_add_35007_comb;
  wire [28:0] p2_add_35022_comb;
  wire [29:0] p2_add_35024_comb;
  wire [30:0] p2_add_35029_comb;
  wire [29:0] p2_add_35030_comb;
  wire [29:0] p2_add_35033_comb;
  wire [29:0] p2_add_35035_comb;
  wire [29:0] p2_add_34115_comb;
  wire [29:0] p2_add_34203_comb;
  wire [31:0] p2_umul_34600_comb;
  wire [31:0] p2_umul_34601_comb;
  wire [29:0] p2_add_34605_comb;
  wire [31:0] p2_umul_34624_comb;
  wire [31:0] p2_umul_34625_comb;
  wire [29:0] p2_add_34629_comb;
  wire [31:0] p2_umul_34632_comb;
  wire [31:0] p2_umul_34633_comb;
  wire [29:0] p2_add_34637_comb;
  wire [31:0] p2_umul_34656_comb;
  wire [31:0] p2_umul_34657_comb;
  wire [29:0] p2_add_34661_comb;
  wire [23:0] p2_bit_slice_34314_comb;
  wire [23:0] p2_bit_slice_34315_comb;
  wire [23:0] p2_bit_slice_34320_comb;
  wire [23:0] p2_bit_slice_34321_comb;
  wire [23:0] p2_bit_slice_34326_comb;
  wire [23:0] p2_bit_slice_34327_comb;
  wire [23:0] p2_bit_slice_34332_comb;
  wire [23:0] p2_bit_slice_34333_comb;
  wire [23:0] p2_bit_slice_34299_comb;
  wire [23:0] p2_bit_slice_34300_comb;
  wire [23:0] p2_bit_slice_34301_comb;
  wire [23:0] p2_bit_slice_34302_comb;
  wire [31:0] p2_sub_35064_comb;
  wire [31:0] p2_sub_35067_comb;
  wire [31:0] p2_sub_35070_comb;
  wire [31:0] p2_concat_34198_comb;
  wire [31:0] p2_concat_34249_comb;
  wire [31:0] p2_or_34692_comb;
  wire [31:0] p2_umul_34693_comb;
  wire [31:0] p2_umul_34694_comb;
  wire [31:0] p2_umul_34696_comb;
  wire [31:0] p2_or_34710_comb;
  wire [31:0] p2_umul_34711_comb;
  wire [31:0] p2_umul_34712_comb;
  wire [31:0] p2_umul_34714_comb;
  wire [31:0] p2_or_34716_comb;
  wire [31:0] p2_umul_34717_comb;
  wire [31:0] p2_umul_34718_comb;
  wire [31:0] p2_umul_34720_comb;
  wire [31:0] p2_or_34734_comb;
  wire [31:0] p2_umul_34735_comb;
  wire [31:0] p2_umul_34736_comb;
  wire [31:0] p2_umul_34738_comb;
  wire [31:0] p2_sub_34349_comb;
  wire [31:0] p2_sub_34350_comb;
  wire [31:0] p2_sign_ext_34351_comb;
  wire [31:0] p2_sign_ext_34352_comb;
  wire [31:0] p2_sub_34353_comb;
  wire [31:0] p2_sub_34354_comb;
  wire [31:0] p2_sign_ext_34355_comb;
  wire [31:0] p2_sign_ext_34356_comb;
  wire [31:0] p2_sub_34361_comb;
  wire [31:0] p2_sub_34362_comb;
  wire [31:0] p2_sign_ext_34363_comb;
  wire [31:0] p2_sign_ext_34364_comb;
  wire [31:0] p2_sub_34365_comb;
  wire [31:0] p2_sub_34366_comb;
  wire [31:0] p2_sign_ext_34367_comb;
  wire [31:0] p2_sign_ext_34368_comb;
  wire [31:0] p2_sign_ext_34334_comb;
  wire [31:0] p2_sign_ext_34335_comb;
  wire [31:0] p2_sign_ext_34336_comb;
  wire [31:0] p2_sign_ext_34337_comb;
  wire [26:0] p2_add_35108_comb;
  wire [26:0] p2_add_35110_comb;
  wire [26:0] p2_add_35112_comb;
  wire [31:0] p2_sub_35093_comb;
  wire [31:0] p2_sub_35096_comb;
  wire [31:0] p2_sub_35099_comb;
  wire [28:0] p2_add_34242_comb;
  wire [31:0] p2_add_34244_comb;
  wire [31:0] p2_add_34245_comb;
  wire [28:0] p2_add_34306_comb;
  wire [31:0] p2_add_34308_comb;
  wire [31:0] p2_add_34309_comb;
  wire [29:0] p2_add_34754_comb;
  wire [31:0] p2_sub_34755_comb;
  wire [31:0] p2_sub_34756_comb;
  wire [31:0] p2_sub_34757_comb;
  wire [29:0] p2_add_34766_comb;
  wire [31:0] p2_sub_34767_comb;
  wire [31:0] p2_sub_34768_comb;
  wire [31:0] p2_sub_34769_comb;
  wire [29:0] p2_add_34770_comb;
  wire [31:0] p2_sub_34771_comb;
  wire [31:0] p2_sub_34772_comb;
  wire [31:0] p2_sub_34773_comb;
  wire [29:0] p2_add_34782_comb;
  wire [31:0] p2_sub_34783_comb;
  wire [31:0] p2_sub_34784_comb;
  wire [31:0] p2_sub_34785_comb;
  wire [23:0] p2_bit_slice_34411_comb;
  wire [23:0] p2_bit_slice_34412_comb;
  wire [31:0] p2_add_34413_comb;
  wire [23:0] p2_bit_slice_34415_comb;
  wire [23:0] p2_bit_slice_34416_comb;
  wire [31:0] p2_add_34417_comb;
  wire [23:0] p2_bit_slice_34423_comb;
  wire [23:0] p2_bit_slice_34424_comb;
  wire [31:0] p2_add_34425_comb;
  wire [23:0] p2_bit_slice_34427_comb;
  wire [23:0] p2_bit_slice_34428_comb;
  wire [31:0] p2_add_34429_comb;
  wire [28:0] p2_concat_35127_comb;
  wire [18:0] p2_add_35114_comb;
  wire [4:0] p2_bit_slice_35115_comb;
  wire [28:0] p2_concat_35128_comb;
  wire [18:0] p2_add_35117_comb;
  wire [4:0] p2_bit_slice_35118_comb;
  wire [28:0] p2_concat_35129_comb;
  wire [18:0] p2_add_35120_comb;
  wire [4:0] p2_bit_slice_35121_comb;
  wire [28:0] p2_bit_slice_34799_comb;
  wire [28:0] p2_bit_slice_34800_comb;
  wire [28:0] p2_bit_slice_34801_comb;
  wire [28:0] p2_bit_slice_34802_comb;
  wire [28:0] p2_bit_slice_34811_comb;
  wire [28:0] p2_bit_slice_34812_comb;
  wire [28:0] p2_bit_slice_34813_comb;
  wire [28:0] p2_bit_slice_34814_comb;
  wire [28:0] p2_bit_slice_34815_comb;
  wire [28:0] p2_bit_slice_34816_comb;
  wire [28:0] p2_bit_slice_34817_comb;
  wire [28:0] p2_bit_slice_34818_comb;
  wire [28:0] p2_bit_slice_34827_comb;
  wire [28:0] p2_bit_slice_34828_comb;
  wire [28:0] p2_bit_slice_34829_comb;
  wire [28:0] p2_bit_slice_34830_comb;
  wire [31:0] p2_sign_ext_34468_comb;
  wire [31:0] p2_sign_ext_34469_comb;
  wire [31:0] p2_umul_34470_comb;
  wire [31:0] p2_sign_ext_34471_comb;
  wire [31:0] p2_sign_ext_34472_comb;
  wire [31:0] p2_umul_34473_comb;
  wire [31:0] p2_sign_ext_34480_comb;
  wire [31:0] p2_sign_ext_34481_comb;
  wire [31:0] p2_umul_34482_comb;
  wire [31:0] p2_sign_ext_34483_comb;
  wire [31:0] p2_sign_ext_34484_comb;
  wire [31:0] p2_umul_34485_comb;
  wire [24:0] p2_add_34433_comb;
  wire [20:0] p2_add_34435_comb;
  wire [24:0] p2_add_34437_comb;
  wire [20:0] p2_add_34439_comb;
  wire [24:0] p2_add_34441_comb;
  wire [20:0] p2_add_34443_comb;
  wire [24:0] p2_add_34445_comb;
  wire [20:0] p2_add_34447_comb;
  wire [24:0] p2_add_34449_comb;
  wire [29:0] p2_add_34450_comb;
  wire [24:0] p2_add_34451_comb;
  wire [29:0] p2_add_34452_comb;
  wire [24:0] p2_add_34453_comb;
  wire [28:0] p2_add_34454_comb;
  wire [24:0] p2_add_34455_comb;
  wire [28:0] p2_add_34456_comb;
  wire [31:0] p2_sign_ext_35136_comb;
  wire [23:0] p2_bit_slice_35116_comb;
  wire [31:0] p2_sign_ext_35138_comb;
  wire [23:0] p2_bit_slice_35119_comb;
  wire [31:0] p2_sign_ext_35140_comb;
  wire [23:0] p2_bit_slice_35122_comb;
  wire [18:0] p2_add_35142_comb;
  wire [18:0] p2_add_35144_comb;
  wire [18:0] p2_add_35146_comb;
  wire [28:0] p2_add_34338_comb;
  wire [30:0] p2_add_34340_comb;
  wire [28:0] p2_add_34342_comb;
  wire [28:0] p2_add_34401_comb;
  wire [30:0] p2_add_34405_comb;
  wire [28:0] p2_add_34407_comb;
  wire [31:0] p2_sign_ext_34853_comb;
  wire [31:0] p2_sign_ext_34854_comb;
  wire [31:0] p2_sign_ext_34855_comb;
  wire [31:0] p2_sign_ext_34856_comb;
  wire [31:0] p2_sign_ext_34857_comb;
  wire [31:0] p2_sign_ext_34858_comb;
  wire [31:0] p2_sign_ext_34859_comb;
  wire [31:0] p2_sign_ext_34860_comb;
  wire [31:0] p2_sign_ext_34861_comb;
  wire [31:0] p2_sign_ext_34862_comb;
  wire [31:0] p2_sign_ext_34863_comb;
  wire [31:0] p2_sign_ext_34864_comb;
  wire [31:0] p2_sign_ext_34865_comb;
  wire [31:0] p2_sign_ext_34866_comb;
  wire [31:0] p2_sign_ext_34867_comb;
  wire [31:0] p2_sign_ext_34868_comb;
  wire [31:0] p2_add_34517_comb;
  wire [31:0] p2_add_34522_comb;
  wire [31:0] p2_add_34537_comb;
  wire [31:0] p2_add_34542_comb;
  wire [23:0] p2_add_35149_comb;
  wire [23:0] p2_add_35151_comb;
  wire [23:0] p2_add_35153_comb;
  wire [23:0] p2_bit_slice_35154_comb;
  wire [23:0] p2_bit_slice_35155_comb;
  wire [23:0] p2_bit_slice_35156_comb;
  wire [31:0] p2_add_34399_comb;
  wire [31:0] p2_add_34459_comb;
  wire [31:0] p2_add_34908_comb;
  wire [31:0] p2_add_34909_comb;
  wire [31:0] p2_add_34910_comb;
  wire [31:0] p2_add_34911_comb;
  wire [31:0] p2_add_34912_comb;
  wire [31:0] p2_add_34913_comb;
  wire [31:0] p2_add_34914_comb;
  wire [31:0] p2_add_34915_comb;
  wire [31:0] p2_add_34995_comb;
  wire [31:0] p2_add_34996_comb;
  wire [31:0] p2_add_35000_comb;
  wire [31:0] p2_add_35001_comb;
  wire [31:0] p2_add_35005_comb;
  wire [31:0] p2_add_35006_comb;
  wire [31:0] p2_add_35010_comb;
  wire [31:0] p2_add_35011_comb;
  wire [31:0] p2_umul_34608_comb;
  wire [31:0] p2_umul_34609_comb;
  wire [29:0] p2_add_34613_comb;
  wire [31:0] p2_umul_34616_comb;
  wire [31:0] p2_umul_34617_comb;
  wire [29:0] p2_add_34621_comb;
  wire [31:0] p2_umul_34640_comb;
  wire [31:0] p2_umul_34641_comb;
  wire [29:0] p2_add_34645_comb;
  wire [31:0] p2_umul_34648_comb;
  wire [31:0] p2_umul_34649_comb;
  wire [29:0] p2_add_34653_comb;
  wire [29:0] p2_add_34551_comb;
  wire [20:0] p2_add_34553_comb;
  wire [29:0] p2_add_34555_comb;
  wire [20:0] p2_add_34557_comb;
  wire [28:0] p2_add_34559_comb;
  wire [20:0] p2_add_34561_comb;
  wire [28:0] p2_add_34563_comb;
  wire [20:0] p2_add_34565_comb;
  wire [20:0] p2_add_34567_comb;
  wire [20:0] p2_add_34570_comb;
  wire [20:0] p2_add_34573_comb;
  wire [20:0] p2_add_34576_comb;
  wire [20:0] p2_add_34579_comb;
  wire [20:0] p2_add_34582_comb;
  wire [20:0] p2_add_34585_comb;
  wire [20:0] p2_add_34588_comb;
  wire [31:0] p2_sub_34919_comb;
  wire [31:0] p2_sub_34968_comb;
  wire [23:0] p2_add_35163_comb;
  wire [23:0] p2_add_35165_comb;
  wire [23:0] p2_add_35167_comb;
  wire [23:0] p2_add_35173_comb;
  wire [31:0] p2_add_35175_comb;
  wire [23:0] p2_add_35176_comb;
  wire [31:0] p2_add_35178_comb;
  wire [23:0] p2_add_35179_comb;
  wire [31:0] p2_add_35181_comb;
  wire [31:0] p2_sub_34457_comb;
  wire [31:0] p2_sub_34461_comb;
  wire [31:0] p2_sub_34506_comb;
  wire [31:0] p2_sub_34509_comb;
  wire [31:0] p2_sub_34951_comb;
  wire [31:0] p2_sub_34953_comb;
  wire [31:0] p2_sub_34955_comb;
  wire [31:0] p2_sub_34957_comb;
  wire [31:0] p2_sub_35044_comb;
  wire [31:0] p2_sub_35048_comb;
  wire [31:0] p2_sub_35052_comb;
  wire [31:0] p2_sub_35056_comb;
  wire [31:0] p2_or_34698_comb;
  wire [31:0] p2_umul_34699_comb;
  wire [31:0] p2_umul_34700_comb;
  wire [31:0] p2_umul_34702_comb;
  wire [31:0] p2_or_34704_comb;
  wire [31:0] p2_umul_34705_comb;
  wire [31:0] p2_umul_34706_comb;
  wire [31:0] p2_umul_34708_comb;
  wire [31:0] p2_or_34722_comb;
  wire [31:0] p2_umul_34723_comb;
  wire [31:0] p2_umul_34724_comb;
  wire [31:0] p2_umul_34726_comb;
  wire [31:0] p2_or_34728_comb;
  wire [31:0] p2_umul_34729_comb;
  wire [31:0] p2_umul_34730_comb;
  wire [31:0] p2_umul_34732_comb;
  wire [31:0] p2_add_34965_comb;
  wire [24:0] p2_add_34966_comb;
  wire [31:0] p2_add_35017_comb;
  wire [24:0] p2_add_35018_comb;
  wire [31:0] p2_add_35183_comb;
  wire [31:0] p2_concat_35184_comb;
  wire [31:0] p2_add_35185_comb;
  wire [31:0] p2_concat_35186_comb;
  wire [31:0] p2_add_35187_comb;
  wire [31:0] p2_concat_35188_comb;
  wire [31:0] p2_sub_35189_comb;
  wire [31:0] p2_sub_35190_comb;
  wire [31:0] p2_sub_35191_comb;
  wire [31:0] p2_add_35193_comb;
  wire [31:0] p2_add_35195_comb;
  wire [31:0] p2_add_35197_comb;
  wire [31:0] p2_umul_34505_comb;
  wire [31:0] p2_umul_34508_comb;
  wire [31:0] p2_umul_34593_comb;
  wire [31:0] p2_umul_34596_comb;
  wire [31:0] p2_umul_34991_comb;
  wire [31:0] p2_umul_34992_comb;
  wire [31:0] p2_umul_34993_comb;
  wire [31:0] p2_umul_34994_comb;
  wire [31:0] p2_umul_35077_comb;
  wire [31:0] p2_umul_35079_comb;
  wire [31:0] p2_umul_35081_comb;
  wire [31:0] p2_umul_35083_comb;
  wire [29:0] p2_add_34758_comb;
  wire [31:0] p2_sub_34759_comb;
  wire [31:0] p2_sub_34760_comb;
  wire [31:0] p2_sub_34761_comb;
  wire [29:0] p2_add_34762_comb;
  wire [31:0] p2_sub_34763_comb;
  wire [31:0] p2_sub_34764_comb;
  wire [31:0] p2_sub_34765_comb;
  wire [29:0] p2_add_34774_comb;
  wire [31:0] p2_sub_34775_comb;
  wire [31:0] p2_sub_34776_comb;
  wire [31:0] p2_sub_34777_comb;
  wire [29:0] p2_add_34778_comb;
  wire [31:0] p2_sub_34779_comb;
  wire [31:0] p2_sub_34780_comb;
  wire [31:0] p2_sub_34781_comb;
  wire [31:0] p2_sub_34739_comb;
  wire [31:0] p2_sub_34740_comb;
  wire [31:0] p2_sub_34741_comb;
  wire [31:0] p2_sub_34742_comb;
  wire [31:0] p2_sub_34743_comb;
  wire [31:0] p2_sub_34744_comb;
  wire [31:0] p2_sub_34745_comb;
  wire [31:0] p2_sub_34746_comb;
  wire [31:0] p2_umul_35047_comb;
  wire [31:0] p2_umul_35051_comb;
  wire [31:0] p2_umul_35055_comb;
  wire [31:0] p2_add_35198_comb;
  wire [31:0] p2_add_35199_comb;
  wire [31:0] p2_add_35200_comb;
  wire [31:0] p2_add_35201_comb;
  wire [31:0] p2_add_35202_comb;
  wire [31:0] p2_add_35203_comb;
  wire [31:0] p2_sub_35204_comb;
  wire [31:0] p2_sub_35205_comb;
  wire [31:0] p2_sub_35206_comb;
  wire [31:0] p2_sub_35207_comb;
  wire [31:0] p2_sub_35208_comb;
  wire [31:0] p2_sub_35209_comb;
  wire [28:0] p2_bit_slice_34803_comb;
  wire [28:0] p2_bit_slice_34804_comb;
  wire [28:0] p2_bit_slice_34805_comb;
  wire [28:0] p2_bit_slice_34806_comb;
  wire [28:0] p2_bit_slice_34807_comb;
  wire [28:0] p2_bit_slice_34808_comb;
  wire [28:0] p2_bit_slice_34809_comb;
  wire [28:0] p2_bit_slice_34810_comb;
  wire [28:0] p2_bit_slice_34819_comb;
  wire [28:0] p2_bit_slice_34820_comb;
  wire [28:0] p2_bit_slice_34821_comb;
  wire [28:0] p2_bit_slice_34822_comb;
  wire [28:0] p2_bit_slice_34823_comb;
  wire [28:0] p2_bit_slice_34824_comb;
  wire [28:0] p2_bit_slice_34825_comb;
  wire [28:0] p2_bit_slice_34826_comb;
  wire [23:0] p2_bit_slice_34786_comb;
  wire [23:0] p2_bit_slice_34787_comb;
  wire [23:0] p2_bit_slice_34788_comb;
  wire [23:0] p2_bit_slice_34789_comb;
  wire [23:0] p2_bit_slice_34790_comb;
  wire [23:0] p2_bit_slice_34791_comb;
  wire [23:0] p2_bit_slice_34792_comb;
  wire [23:0] p2_bit_slice_34793_comb;
  wire [29:0] p2_add_35061_comb;
  wire [31:0] p2_sub_35078_comb;
  wire [31:0] p2_sub_35080_comb;
  wire [31:0] p2_sub_35082_comb;
  wire [29:0] p2_add_35090_comb;
  wire [31:0] p2_add_35172_comb;
  wire [31:0] p2_add_35182_comb;
  wire [17:0] p2_bit_slice_35210_comb;
  wire [17:0] p2_bit_slice_35211_comb;
  wire [17:0] p2_bit_slice_35212_comb;
  wire [17:0] p2_bit_slice_35213_comb;
  wire [17:0] p2_bit_slice_35214_comb;
  wire [17:0] p2_bit_slice_35215_comb;
  wire [17:0] p2_bit_slice_35216_comb;
  wire [17:0] p2_bit_slice_35217_comb;
  wire [17:0] p2_bit_slice_35218_comb;
  wire [17:0] p2_bit_slice_35219_comb;
  wire [17:0] p2_bit_slice_35220_comb;
  wire [17:0] p2_bit_slice_35221_comb;
  wire [24:0] p2_add_34680_comb;
  wire [24:0] p2_add_34683_comb;
  wire [24:0] p2_add_34747_comb;
  wire [24:0] p2_add_34749_comb;
  wire [24:0] p2_add_35073_comb;
  wire [24:0] p2_add_35074_comb;
  wire [24:0] p2_add_35075_comb;
  wire [24:0] p2_add_35076_comb;
  wire [24:0] p2_add_35123_comb;
  wire [24:0] p2_add_35124_comb;
  wire [24:0] p2_add_35125_comb;
  wire [24:0] p2_add_35126_comb;
  wire [31:0] p2_umul_34794_comb;
  wire [31:0] p2_umul_34837_comb;
  assign p2_umul_33941_comb = umul32b_32b_x_8b(p1_sub_33085, 8'hb5);
  assign p2_umul_33942_comb = umul32b_32b_x_8b(p1_sub_33086, 8'hb5);
  assign p2_umul_33943_comb = umul32b_32b_x_8b(p1_sub_33095, 8'hb5);
  assign p2_umul_33944_comb = umul32b_32b_x_8b(p1_sub_33096, 8'hb5);
  assign p2_umul_33957_comb = umul32b_32b_x_8b(p1_sub_33135, 8'hb5);
  assign p2_umul_33958_comb = umul32b_32b_x_8b(p1_sub_33136, 8'hb5);
  assign p2_add_33959_comb = p2_umul_33941_comb[31:7] + 25'h000_0001;
  assign p2_add_33960_comb = p2_umul_33942_comb[31:7] + 25'h000_0001;
  assign p2_umul_33961_comb = umul32b_32b_x_8b(p1_sub_33137, 8'hb5);
  assign p2_umul_33962_comb = umul32b_32b_x_8b(p1_sub_33138, 8'hb5);
  assign p2_add_33963_comb = p2_umul_33943_comb[31:7] + 25'h000_0001;
  assign p2_add_33964_comb = p2_umul_33944_comb[31:7] + 25'h000_0001;
  assign p2_add_34598_comb = p1_array_index_33709 + p1_array_index_33710;
  assign p2_bit_slice_33969_comb = p2_add_33959_comb[24:1];
  assign p2_bit_slice_33970_comb = p2_add_33960_comb[24:1];
  assign p2_bit_slice_33975_comb = p2_add_33963_comb[24:1];
  assign p2_bit_slice_33976_comb = p2_add_33964_comb[24:1];
  assign p2_umul_34686_comb = umul32b_32b_x_11b(p1_array_index_33709, 11'h620);
  assign p2_umul_34687_comb = umul32b_32b_x_11b(p2_add_34598_comb, 11'h454);
  assign p2_add_34689_comb = p1_array_index_33739 + p1_array_index_33740;
  assign p2_add_33977_comb = p2_umul_33957_comb[31:7] + 25'h000_0001;
  assign p2_add_33978_comb = p2_umul_33958_comb[31:7] + 25'h000_0001;
  assign p2_sign_ext_33979_comb = {{8{p2_bit_slice_33969_comb[23]}}, p2_bit_slice_33969_comb};
  assign p2_sign_ext_33980_comb = {{8{p2_bit_slice_33970_comb[23]}}, p2_bit_slice_33970_comb};
  assign p2_add_33981_comb = p2_umul_33961_comb[31:7] + 25'h000_0001;
  assign p2_add_33982_comb = p2_umul_33962_comb[31:7] + 25'h000_0001;
  assign p2_sign_ext_33983_comb = {{8{p2_bit_slice_33975_comb[23]}}, p2_bit_slice_33975_comb};
  assign p2_sign_ext_33984_comb = {{8{p2_bit_slice_33976_comb[23]}}, p2_bit_slice_33976_comb};
  assign p2_add_34057_comb = p1_array_index_33285 + p1_array_index_33286;
  assign p2_add_33986_comb = p1_array_index_33203 + p1_array_index_33204;
  assign p2_umul_34752_comb = umul32b_32b_x_11b(p1_array_index_33739, 11'h620);
  assign p2_umul_34753_comb = umul32b_32b_x_11b(p2_add_34689_comb, 11'h454);
  assign p2_bit_slice_33988_comb = p2_add_33977_comb[24:1];
  assign p2_bit_slice_33989_comb = p2_add_33978_comb[24:1];
  assign p2_bit_slice_33996_comb = p2_add_33981_comb[24:1];
  assign p2_bit_slice_33997_comb = p2_add_33982_comb[24:1];
  assign p2_umul_34112_comb = umul32b_32b_x_12b(p2_add_34057_comb, 12'h968);
  assign p2_umul_34021_comb = umul32b_32b_x_10b(p2_add_33986_comb, 10'h235);
  assign p2_umul_34199_comb = umul32b_32b_x_12b(p1_array_index_33286, 12'hfb1);
  assign p2_umul_34113_comb = umul32b_32b_x_12b(p1_array_index_33204, 12'hd4e);
  assign p2_umul_34197_comb = umul32b_32b_x_10b(p1_array_index_33285, 10'h31f);
  assign p2_add_34796_comb = p2_umul_34686_comb[31:5] + p2_umul_34687_comb[31:5];
  assign p2_umul_34020_comb = umul32b_32b_x_12b(p1_array_index_33203, 12'h8e4);
  assign p2_add_34118_comb = p1_array_index_33343 + p1_array_index_33344;
  assign p2_add_34023_comb = p1_array_index_33237 + p1_array_index_33238;
  assign p2_sign_ext_34025_comb = {{8{p2_bit_slice_33988_comb[23]}}, p2_bit_slice_33988_comb};
  assign p2_sign_ext_34026_comb = {{8{p2_bit_slice_33989_comb[23]}}, p2_bit_slice_33989_comb};
  assign p2_add_34027_comb = p2_sign_ext_33979_comb[31:7] + 25'h000_0001;
  assign p2_add_34029_comb = p1_umul_33168[31:11] + p1_bit_slice_33214;
  assign p2_add_34031_comb = p2_sign_ext_33980_comb[31:7] + 25'h000_0001;
  assign p2_add_34033_comb = p1_umul_33170[31:11] + p1_bit_slice_33216;
  assign p2_sign_ext_34035_comb = {{8{p2_bit_slice_33996_comb[23]}}, p2_bit_slice_33996_comb};
  assign p2_sign_ext_34036_comb = {{8{p2_bit_slice_33997_comb[23]}}, p2_bit_slice_33997_comb};
  assign p2_add_34037_comb = p2_sign_ext_33983_comb[31:7] + 25'h000_0001;
  assign p2_add_34039_comb = p1_umul_33207[31:11] + p1_bit_slice_33214;
  assign p2_add_34041_comb = p2_sign_ext_33984_comb[31:7] + 25'h000_0001;
  assign p2_add_34043_comb = p1_umul_33208[31:11] + p1_bit_slice_33216;
  assign p2_add_34045_comb = p1_umul_33207[31:7] + 25'h000_0001;
  assign p2_add_34046_comb = p2_sign_ext_33983_comb[31:2] + p1_umul_33168[31:2];
  assign p2_add_34047_comb = p1_umul_33208[31:7] + 25'h000_0001;
  assign p2_add_34048_comb = p2_sign_ext_33984_comb[31:2] + p1_umul_33170[31:2];
  assign p2_add_34049_comb = p1_umul_33168[31:7] + 25'h000_0001;
  assign p2_add_34050_comb = p2_sign_ext_33979_comb[31:3] + p1_umul_33207[31:3];
  assign p2_add_34051_comb = p1_umul_33170[31:7] + 25'h000_0001;
  assign p2_add_34052_comb = p2_sign_ext_33980_comb[31:3] + p1_umul_33208[31:3];
  assign p2_sign_ext_34831_comb = {{8{p1_bit_slice_33773[23]}}, p1_bit_slice_33773};
  assign p2_sign_ext_34832_comb = {{8{p1_bit_slice_33774[23]}}, p1_bit_slice_33774};
  assign p2_add_34841_comb = p1_bit_slice_33779 + p1_bit_slice_33780;
  assign p2_sign_ext_34833_comb = {{8{p1_bit_slice_33775[23]}}, p1_bit_slice_33775};
  assign p2_sign_ext_34834_comb = {{8{p1_bit_slice_33776[23]}}, p1_bit_slice_33776};
  assign p2_sign_ext_34835_comb = {{8{p1_bit_slice_33777[23]}}, p1_bit_slice_33777};
  assign p2_sign_ext_34836_comb = {{8{p1_bit_slice_33778[23]}}, p1_bit_slice_33778};
  assign p2_umul_34200_comb = umul32b_32b_x_12b(p2_add_34118_comb, 12'h968);
  assign p2_umul_34063_comb = umul32b_32b_x_10b(p2_add_34023_comb, 10'h235);
  assign p2_umul_34250_comb = umul32b_32b_x_12b(p1_array_index_33344, 12'hfb1);
  assign p2_umul_34201_comb = umul32b_32b_x_12b(p1_array_index_33238, 12'hd4e);
  assign p2_umul_34248_comb = umul32b_32b_x_10b(p1_array_index_33343, 10'h31f);
  assign p2_add_34852_comb = p2_umul_34752_comb[31:5] + p2_umul_34753_comb[31:5];
  assign p2_umul_34062_comb = umul32b_32b_x_12b(p1_array_index_33237, 12'h8e4);
  assign p2_sign_ext_34347_comb = {{8{p1_bit_slice_33571[23]}}, p1_bit_slice_33571};
  assign p2_sign_ext_34348_comb = {{8{p1_bit_slice_33572[23]}}, p1_bit_slice_33572};
  assign p2_sign_ext_34357_comb = {{8{p1_bit_slice_33577[23]}}, p1_bit_slice_33577};
  assign p2_sign_ext_34358_comb = {{8{p1_bit_slice_33578[23]}}, p1_bit_slice_33578};
  assign p2_sign_ext_34359_comb = {{8{p1_bit_slice_33583[23]}}, p1_bit_slice_33583};
  assign p2_sign_ext_34360_comb = {{8{p1_bit_slice_33584[23]}}, p1_bit_slice_33584};
  assign p2_sign_ext_34369_comb = {{8{p1_bit_slice_33589[23]}}, p1_bit_slice_33589};
  assign p2_sign_ext_34370_comb = {{8{p1_bit_slice_33590[23]}}, p1_bit_slice_33590};
  assign p2_add_34869_comb = p2_sign_ext_34831_comb + p2_sign_ext_34832_comb;
  assign p2_add_34876_comb = p2_umul_34112_comb[31:7] + 25'h000_0001;
  assign p2_add_34878_comb = p2_umul_34021_comb[31:11] + p2_add_34841_comb;
  assign p2_add_34880_comb = p2_umul_34199_comb[31:1] + p2_umul_34113_comb[31:1];
  assign p2_add_34871_comb = p2_sign_ext_34833_comb + p2_sign_ext_34834_comb;
  assign p2_add_34888_comb = p2_umul_34199_comb[31:7] + 25'h000_0001;
  assign p2_add_34890_comb = p2_umul_34113_comb[31:11] + p2_add_34841_comb;
  assign p2_add_34892_comb = p2_umul_34112_comb[31:3] + p2_umul_34021_comb[31:3];
  assign p2_add_34873_comb = p2_sign_ext_34835_comb + p2_sign_ext_34836_comb;
  assign p2_add_34898_comb = p2_umul_34197_comb[31:7] + 25'h000_0001;
  assign p2_add_34900_comb = p2_add_34796_comb[26:6] + p2_add_34841_comb;
  assign p2_add_34902_comb = p2_umul_34112_comb[31:3] + p2_umul_34020_comb[31:3];
  assign p2_add_34885_comb = p1_bit_slice_33783 + p1_bit_slice_33784;
  assign p2_add_34409_comb = p2_sign_ext_34347_comb + p2_sign_ext_34348_comb;
  assign p2_add_34419_comb = p2_sign_ext_34357_comb + p2_sign_ext_34358_comb;
  assign p2_add_34421_comb = p2_sign_ext_34359_comb + p2_sign_ext_34360_comb;
  assign p2_add_34431_comb = p2_sign_ext_34369_comb + p2_sign_ext_34370_comb;
  assign p2_add_34123_comb = p2_sign_ext_34025_comb[31:7] + 25'h000_0001;
  assign p2_add_34125_comb = p1_umul_33218[31:11] + p1_bit_slice_33294;
  assign p2_add_34127_comb = p2_sign_ext_34026_comb[31:7] + 25'h000_0001;
  assign p2_add_34129_comb = p1_umul_33220[31:11] + p1_bit_slice_33296;
  assign p2_add_34131_comb = {p2_add_34027_comb, p2_add_33959_comb[7:3]} + {p2_add_34029_comb, p1_umul_33168[10:2]};
  assign p2_add_34133_comb = p1_umul_33207[31:11] + p1_bit_slice_33213;
  assign p2_add_34135_comb = {p2_add_34031_comb, p2_add_33960_comb[7:3]} + {p2_add_34033_comb, p1_umul_33170[10:2]};
  assign p2_add_34137_comb = p1_umul_33208[31:11] + p1_bit_slice_33215;
  assign p2_add_34139_comb = p2_sign_ext_34035_comb[31:7] + 25'h000_0001;
  assign p2_add_34141_comb = p1_umul_33291[31:11] + p1_bit_slice_33294;
  assign p2_add_34143_comb = p2_sign_ext_34036_comb[31:7] + 25'h000_0001;
  assign p2_add_34145_comb = p1_umul_33292[31:11] + p1_bit_slice_33296;
  assign p2_add_34147_comb = {p2_add_34037_comb, p2_add_33963_comb[7:4]} + {p2_add_34039_comb, p1_umul_33207[10:3]};
  assign p2_add_34149_comb = p1_umul_33168[31:11] + p1_bit_slice_33213;
  assign p2_add_34151_comb = {p2_add_34041_comb, p2_add_33964_comb[7:4]} + {p2_add_34043_comb, p1_umul_33208[10:3]};
  assign p2_add_34153_comb = p1_umul_33170[31:11] + p1_bit_slice_33215;
  assign p2_add_34155_comb = p1_umul_33291[31:7] + 25'h000_0001;
  assign p2_add_34156_comb = p2_sign_ext_34035_comb[31:2] + p1_umul_33218[31:2];
  assign p2_add_34157_comb = p1_umul_33292[31:7] + 25'h000_0001;
  assign p2_add_34158_comb = p2_sign_ext_34036_comb[31:2] + p1_umul_33220[31:2];
  assign p2_add_34159_comb = p2_add_34045_comb[24:4] + p1_bit_slice_33214;
  assign p2_add_34162_comb = p2_add_34046_comb[29:9] + p1_bit_slice_33213;
  assign p2_add_34165_comb = p2_add_34047_comb[24:4] + p1_bit_slice_33216;
  assign p2_add_34168_comb = p2_add_34048_comb[29:9] + p1_bit_slice_33215;
  assign p2_add_34171_comb = p1_umul_33218[31:7] + 25'h000_0001;
  assign p2_add_34172_comb = p2_sign_ext_34025_comb[31:3] + p1_umul_33291[31:3];
  assign p2_add_34173_comb = p1_umul_33220[31:7] + 25'h000_0001;
  assign p2_add_34174_comb = p2_sign_ext_34026_comb[31:3] + p1_umul_33292[31:3];
  assign p2_add_34175_comb = p2_add_34049_comb[24:4] + p1_bit_slice_33214;
  assign p2_add_34178_comb = p2_add_34050_comb[28:8] + p1_bit_slice_33213;
  assign p2_add_34181_comb = p2_add_34051_comb[24:4] + p1_bit_slice_33216;
  assign p2_add_34184_comb = p2_add_34052_comb[28:8] + p1_bit_slice_33215;
  assign p2_umul_34108_comb = umul32b_32b_x_8b(p1_sub_33335, 8'hb5);
  assign p2_umul_34109_comb = umul32b_32b_x_8b(p1_sub_33336, 8'hb5);
  assign p2_umul_34110_comb = umul32b_32b_x_8b(p1_sub_33337, 8'hb5);
  assign p2_umul_34111_comb = umul32b_32b_x_8b(p1_sub_33338, 8'hb5);
  assign p2_umul_34916_comb = umul32b_32b_x_11b(p2_add_34869_comb, 11'h454);
  assign p2_concat_34926_comb = {p2_add_34796_comb, p2_umul_34687_comb[4:2]};
  assign p2_umul_34917_comb = umul32b_32b_x_11b(p2_add_34871_comb, 11'h454);
  assign p2_umul_34918_comb = umul32b_32b_x_11b(p2_add_34873_comb, 11'h454);
  assign p2_add_34927_comb = p2_umul_34200_comb[31:7] + 25'h000_0001;
  assign p2_add_34929_comb = p2_umul_34063_comb[31:11] + p2_add_34885_comb;
  assign p2_add_34931_comb = p2_umul_34250_comb[31:1] + p2_umul_34201_comb[31:1];
  assign p2_add_34936_comb = p2_umul_34250_comb[31:7] + 25'h000_0001;
  assign p2_add_34938_comb = p2_umul_34201_comb[31:11] + p2_add_34885_comb;
  assign p2_add_34940_comb = p2_umul_34200_comb[31:3] + p2_umul_34063_comb[31:3];
  assign p2_add_34945_comb = p2_umul_34248_comb[31:7] + 25'h000_0001;
  assign p2_add_34947_comb = p2_add_34852_comb[26:6] + p2_add_34885_comb;
  assign p2_add_34949_comb = p2_umul_34200_comb[31:3] + p2_umul_34062_comb[31:3];
  assign p2_sign_ext_34465_comb = {{8{p1_bit_slice_33635[23]}}, p1_bit_slice_33635};
  assign p2_sign_ext_34466_comb = {{8{p1_bit_slice_33636[23]}}, p1_bit_slice_33636};
  assign p2_umul_34467_comb = umul32b_32b_x_10b(p2_add_34409_comb, 10'h235);
  assign p2_sign_ext_34474_comb = {{8{p1_bit_slice_33637[23]}}, p1_bit_slice_33637};
  assign p2_sign_ext_34475_comb = {{8{p1_bit_slice_33638[23]}}, p1_bit_slice_33638};
  assign p2_umul_34476_comb = umul32b_32b_x_10b(p2_add_34419_comb, 10'h235);
  assign p2_sign_ext_34477_comb = {{8{p1_bit_slice_33639[23]}}, p1_bit_slice_33639};
  assign p2_sign_ext_34478_comb = {{8{p1_bit_slice_33640[23]}}, p1_bit_slice_33640};
  assign p2_umul_34479_comb = umul32b_32b_x_10b(p2_add_34421_comb, 10'h235);
  assign p2_sign_ext_34486_comb = {{8{p1_bit_slice_33641[23]}}, p1_bit_slice_33641};
  assign p2_sign_ext_34487_comb = {{8{p1_bit_slice_33642[23]}}, p1_bit_slice_33642};
  assign p2_umul_34488_comb = umul32b_32b_x_10b(p2_add_34431_comb, 10'h235);
  assign p2_add_34971_comb = {p2_add_34876_comb, p2_umul_34112_comb[6:3]} + {p2_add_34878_comb, p2_umul_34021_comb[10:3]};
  assign p2_add_34973_comb = p2_add_34880_comb[30:1] + p2_concat_34926_comb;
  assign p2_add_34980_comb = {p2_add_34888_comb, p2_umul_34199_comb[6:1]} + {p2_add_34890_comb, p2_umul_34113_comb[10:1]};
  assign p2_add_34981_comb = {p2_add_34892_comb, p2_umul_34021_comb[2]} + p2_concat_34926_comb;
  assign p2_add_34985_comb = {p2_add_34898_comb, p2_umul_34197_comb[6:2]} + {p2_add_34900_comb, p2_add_34796_comb[5:0], p2_umul_34687_comb[4:2]};
  assign p2_add_34987_comb = {p2_add_34902_comb, p2_umul_34020_comb[2]} + p2_umul_34021_comb[31:2];
  assign p2_concat_34979_comb = {p2_add_34852_comb, p2_umul_34753_comb[4:2]};
  assign p2_add_34512_comb = p2_sign_ext_34465_comb + p2_sign_ext_34466_comb;
  assign p2_add_34527_comb = p2_sign_ext_34474_comb + p2_sign_ext_34475_comb;
  assign p2_add_34532_comb = p2_sign_ext_34477_comb + p2_sign_ext_34478_comb;
  assign p2_add_34547_comb = p2_sign_ext_34486_comb + p2_sign_ext_34487_comb;
  assign p2_add_34251_comb = {p2_add_34123_comb, p2_add_33977_comb[7:3]} + {p2_add_34125_comb, p1_umul_33218[10:2]};
  assign p2_add_34253_comb = p1_umul_33291[31:11] + p1_bit_slice_33293;
  assign p2_add_34255_comb = {p2_add_34127_comb, p2_add_33978_comb[7:3]} + {p2_add_34129_comb, p1_umul_33220[10:2]};
  assign p2_add_34257_comb = p1_umul_33292[31:11] + p1_bit_slice_33295;
  assign p2_sub_34259_comb = {p2_add_34131_comb, p2_add_33959_comb[2:1]} - {p2_add_34133_comb, p1_umul_33207[10:0]};
  assign p2_sub_34260_comb = {p2_add_34135_comb, p2_add_33960_comb[2:1]} - {p2_add_34137_comb, p1_umul_33208[10:0]};
  assign p2_add_34261_comb = {p2_add_34139_comb, p2_add_33981_comb[7:4]} + {p2_add_34141_comb, p1_umul_33291[10:3]};
  assign p2_add_34263_comb = p1_umul_33218[31:11] + p1_bit_slice_33293;
  assign p2_add_34265_comb = {p2_add_34143_comb, p2_add_33982_comb[7:4]} + {p2_add_34145_comb, p1_umul_33292[10:3]};
  assign p2_add_34267_comb = p1_umul_33220[31:11] + p1_bit_slice_33295;
  assign p2_sub_34269_comb = {p2_add_34147_comb, p2_add_33963_comb[3:1]} - {p2_add_34149_comb, p1_umul_33168[10:0]};
  assign p2_sub_34270_comb = {p2_add_34151_comb, p2_add_33964_comb[3:1]} - {p2_add_34153_comb, p1_umul_33170[10:0]};
  assign p2_add_34271_comb = p2_add_34155_comb[24:4] + p1_bit_slice_33294;
  assign p2_add_34274_comb = p2_add_34156_comb[29:9] + p1_bit_slice_33293;
  assign p2_add_34277_comb = p2_add_34157_comb[24:4] + p1_bit_slice_33296;
  assign p2_add_34280_comb = p2_add_34158_comb[29:9] + p1_bit_slice_33295;
  assign p2_sub_34283_comb = {p2_add_34159_comb, p2_add_34045_comb[3:0], p1_umul_33207[6:0]} - {p2_add_34162_comb, p2_add_34046_comb[8:0], p2_add_33963_comb[2:1]};
  assign p2_sub_34284_comb = {p2_add_34165_comb, p2_add_34047_comb[3:0], p1_umul_33208[6:0]} - {p2_add_34168_comb, p2_add_34048_comb[8:0], p2_add_33964_comb[2:1]};
  assign p2_add_34285_comb = p2_add_34171_comb[24:4] + p1_bit_slice_33294;
  assign p2_add_34288_comb = p2_add_34172_comb[28:8] + p1_bit_slice_33293;
  assign p2_add_34291_comb = p2_add_34173_comb[24:4] + p1_bit_slice_33296;
  assign p2_add_34294_comb = p2_add_34174_comb[28:8] + p1_bit_slice_33295;
  assign p2_sub_34297_comb = {p2_add_34175_comb, p2_add_34049_comb[3:0], p1_umul_33168[6:0]} - {p2_add_34178_comb, p2_add_34050_comb[7:0], p2_add_33959_comb[3:1]};
  assign p2_sub_34298_comb = {p2_add_34181_comb, p2_add_34051_comb[3:0], p1_umul_33170[6:0]} - {p2_add_34184_comb, p2_add_34052_comb[7:0], p2_add_33960_comb[3:1]};
  assign p2_add_34238_comb = p2_umul_34108_comb[31:7] + 25'h000_0001;
  assign p2_add_34239_comb = p2_umul_34109_comb[31:7] + 25'h000_0001;
  assign p2_add_34240_comb = p2_umul_34110_comb[31:7] + 25'h000_0001;
  assign p2_add_34241_comb = p2_umul_34111_comb[31:7] + 25'h000_0001;
  assign p2_umul_35058_comb = umul32b_32b_x_11b(p2_sign_ext_34831_comb, 11'h620);
  assign p2_add_34997_comb = p2_umul_34916_comb[31:2] + 30'h0000_0001;
  assign p2_umul_35059_comb = umul32b_32b_x_11b(p2_sign_ext_34833_comb, 11'h620);
  assign p2_add_35002_comb = p2_umul_34917_comb[31:2] + 30'h0000_0001;
  assign p2_umul_35060_comb = umul32b_32b_x_11b(p2_sign_ext_34835_comb, 11'h620);
  assign p2_add_35007_comb = p2_umul_34918_comb[31:2] + 30'h0000_0001;
  assign p2_add_35022_comb = {p2_add_34927_comb, p2_umul_34200_comb[6:3]} + {p2_add_34929_comb, p2_umul_34063_comb[10:3]};
  assign p2_add_35024_comb = p2_add_34931_comb[30:1] + p2_concat_34979_comb;
  assign p2_add_35029_comb = {p2_add_34936_comb, p2_umul_34250_comb[6:1]} + {p2_add_34938_comb, p2_umul_34201_comb[10:1]};
  assign p2_add_35030_comb = {p2_add_34940_comb, p2_umul_34063_comb[2]} + p2_concat_34979_comb;
  assign p2_add_35033_comb = {p2_add_34945_comb, p2_umul_34248_comb[6:2]} + {p2_add_34947_comb, p2_add_34852_comb[5:0], p2_umul_34753_comb[4:2]};
  assign p2_add_35035_comb = {p2_add_34949_comb, p2_umul_34062_comb[2]} + p2_umul_34063_comb[31:2];
  assign p2_add_34115_comb = p2_umul_34020_comb[31:2] + p2_umul_34021_comb[31:2];
  assign p2_add_34203_comb = p2_umul_34062_comb[31:2] + p2_umul_34063_comb[31:2];
  assign p2_umul_34600_comb = umul32b_32b_x_12b(p2_sign_ext_34347_comb, 12'h8e4);
  assign p2_umul_34601_comb = umul32b_32b_x_12b(p2_add_34512_comb, 12'h968);
  assign p2_add_34605_comb = p2_umul_34467_comb[31:2] + 30'h0000_0001;
  assign p2_umul_34624_comb = umul32b_32b_x_12b(p2_sign_ext_34357_comb, 12'h8e4);
  assign p2_umul_34625_comb = umul32b_32b_x_12b(p2_add_34527_comb, 12'h968);
  assign p2_add_34629_comb = p2_umul_34476_comb[31:2] + 30'h0000_0001;
  assign p2_umul_34632_comb = umul32b_32b_x_12b(p2_sign_ext_34359_comb, 12'h8e4);
  assign p2_umul_34633_comb = umul32b_32b_x_12b(p2_add_34532_comb, 12'h968);
  assign p2_add_34637_comb = p2_umul_34479_comb[31:2] + 30'h0000_0001;
  assign p2_umul_34656_comb = umul32b_32b_x_12b(p2_sign_ext_34369_comb, 12'h8e4);
  assign p2_umul_34657_comb = umul32b_32b_x_12b(p2_add_34547_comb, 12'h968);
  assign p2_add_34661_comb = p2_umul_34488_comb[31:2] + 30'h0000_0001;
  assign p2_bit_slice_34314_comb = p2_sub_34259_comb[31:8];
  assign p2_bit_slice_34315_comb = p2_sub_34260_comb[31:8];
  assign p2_bit_slice_34320_comb = p2_sub_34269_comb[31:8];
  assign p2_bit_slice_34321_comb = p2_sub_34270_comb[31:8];
  assign p2_bit_slice_34326_comb = p2_sub_34283_comb[31:8];
  assign p2_bit_slice_34327_comb = p2_sub_34284_comb[31:8];
  assign p2_bit_slice_34332_comb = p2_sub_34297_comb[31:8];
  assign p2_bit_slice_34333_comb = p2_sub_34298_comb[31:8];
  assign p2_bit_slice_34299_comb = p2_add_34238_comb[24:1];
  assign p2_bit_slice_34300_comb = p2_add_34239_comb[24:1];
  assign p2_bit_slice_34301_comb = p2_add_34240_comb[24:1];
  assign p2_bit_slice_34302_comb = p2_add_34241_comb[24:1];
  assign p2_sub_35064_comb = {p2_add_34971_comb, p2_umul_34021_comb[2:0]} - {p2_add_34973_comb, p2_add_34880_comb[0], p2_umul_34199_comb[0]};
  assign p2_sub_35067_comb = {p2_add_34980_comb, p2_umul_34199_comb[0]} - {p2_add_34981_comb, p2_umul_34021_comb[1:0]};
  assign p2_sub_35070_comb = {p2_add_34985_comb, p2_umul_34197_comb[1:0]} - {p2_add_34987_comb, p2_umul_34021_comb[1:0]};
  assign p2_concat_34198_comb = {p2_add_34115_comb, p2_umul_34021_comb[1:0]};
  assign p2_concat_34249_comb = {p2_add_34203_comb, p2_umul_34063_comb[1:0]};
  assign p2_or_34692_comb = p2_umul_34601_comb | 32'h0000_0004;
  assign p2_umul_34693_comb = umul32b_32b_x_12b(p2_sign_ext_34466_comb, 12'hfb1);
  assign p2_umul_34694_comb = umul32b_32b_x_10b(p2_sign_ext_34465_comb, 10'h31f);
  assign p2_umul_34696_comb = umul32b_32b_x_12b(p2_sign_ext_34348_comb, 12'hd4e);
  assign p2_or_34710_comb = p2_umul_34625_comb | 32'h0000_0004;
  assign p2_umul_34711_comb = umul32b_32b_x_12b(p2_sign_ext_34475_comb, 12'hfb1);
  assign p2_umul_34712_comb = umul32b_32b_x_10b(p2_sign_ext_34474_comb, 10'h31f);
  assign p2_umul_34714_comb = umul32b_32b_x_12b(p2_sign_ext_34358_comb, 12'hd4e);
  assign p2_or_34716_comb = p2_umul_34633_comb | 32'h0000_0004;
  assign p2_umul_34717_comb = umul32b_32b_x_12b(p2_sign_ext_34478_comb, 12'hfb1);
  assign p2_umul_34718_comb = umul32b_32b_x_10b(p2_sign_ext_34477_comb, 10'h31f);
  assign p2_umul_34720_comb = umul32b_32b_x_12b(p2_sign_ext_34360_comb, 12'hd4e);
  assign p2_or_34734_comb = p2_umul_34657_comb | 32'h0000_0004;
  assign p2_umul_34735_comb = umul32b_32b_x_12b(p2_sign_ext_34487_comb, 12'hfb1);
  assign p2_umul_34736_comb = umul32b_32b_x_10b(p2_sign_ext_34486_comb, 10'h31f);
  assign p2_umul_34738_comb = umul32b_32b_x_12b(p2_sign_ext_34370_comb, 12'hd4e);
  assign p2_sub_34349_comb = {p2_add_34251_comb, p2_add_33977_comb[2:1]} - {p2_add_34253_comb, p1_umul_33291[10:0]};
  assign p2_sub_34350_comb = {p2_add_34255_comb, p2_add_33978_comb[2:1]} - {p2_add_34257_comb, p1_umul_33292[10:0]};
  assign p2_sign_ext_34351_comb = {{8{p2_bit_slice_34314_comb[23]}}, p2_bit_slice_34314_comb};
  assign p2_sign_ext_34352_comb = {{8{p2_bit_slice_34315_comb[23]}}, p2_bit_slice_34315_comb};
  assign p2_sub_34353_comb = {p2_add_34261_comb, p2_add_33981_comb[3:1]} - {p2_add_34263_comb, p1_umul_33218[10:0]};
  assign p2_sub_34354_comb = {p2_add_34265_comb, p2_add_33982_comb[3:1]} - {p2_add_34267_comb, p1_umul_33220[10:0]};
  assign p2_sign_ext_34355_comb = {{8{p2_bit_slice_34320_comb[23]}}, p2_bit_slice_34320_comb};
  assign p2_sign_ext_34356_comb = {{8{p2_bit_slice_34321_comb[23]}}, p2_bit_slice_34321_comb};
  assign p2_sub_34361_comb = {p2_add_34271_comb, p2_add_34155_comb[3:0], p1_umul_33291[6:0]} - {p2_add_34274_comb, p2_add_34156_comb[8:0], p2_add_33981_comb[2:1]};
  assign p2_sub_34362_comb = {p2_add_34277_comb, p2_add_34157_comb[3:0], p1_umul_33292[6:0]} - {p2_add_34280_comb, p2_add_34158_comb[8:0], p2_add_33982_comb[2:1]};
  assign p2_sign_ext_34363_comb = {{8{p2_bit_slice_34326_comb[23]}}, p2_bit_slice_34326_comb};
  assign p2_sign_ext_34364_comb = {{8{p2_bit_slice_34327_comb[23]}}, p2_bit_slice_34327_comb};
  assign p2_sub_34365_comb = {p2_add_34285_comb, p2_add_34171_comb[3:0], p1_umul_33218[6:0]} - {p2_add_34288_comb, p2_add_34172_comb[7:0], p2_add_33977_comb[3:1]};
  assign p2_sub_34366_comb = {p2_add_34291_comb, p2_add_34173_comb[3:0], p1_umul_33220[6:0]} - {p2_add_34294_comb, p2_add_34174_comb[7:0], p2_add_33978_comb[3:1]};
  assign p2_sign_ext_34367_comb = {{8{p2_bit_slice_34332_comb[23]}}, p2_bit_slice_34332_comb};
  assign p2_sign_ext_34368_comb = {{8{p2_bit_slice_34333_comb[23]}}, p2_bit_slice_34333_comb};
  assign p2_sign_ext_34334_comb = {{8{p2_bit_slice_34299_comb[23]}}, p2_bit_slice_34299_comb};
  assign p2_sign_ext_34335_comb = {{8{p2_bit_slice_34300_comb[23]}}, p2_bit_slice_34300_comb};
  assign p2_sign_ext_34336_comb = {{8{p2_bit_slice_34301_comb[23]}}, p2_bit_slice_34301_comb};
  assign p2_sign_ext_34337_comb = {{8{p2_bit_slice_34302_comb[23]}}, p2_bit_slice_34302_comb};
  assign p2_add_35108_comb = p2_umul_35058_comb[31:5] + p2_add_34997_comb[29:3];
  assign p2_add_35110_comb = p2_umul_35059_comb[31:5] + p2_add_35002_comb[29:3];
  assign p2_add_35112_comb = p2_umul_35060_comb[31:5] + p2_add_35007_comb[29:3];
  assign p2_sub_35093_comb = {p2_add_35022_comb, p2_umul_34063_comb[2:0]} - {p2_add_35024_comb, p2_add_34931_comb[0], p2_umul_34250_comb[0]};
  assign p2_sub_35096_comb = {p2_add_35029_comb, p2_umul_34250_comb[0]} - {p2_add_35030_comb, p2_umul_34063_comb[1:0]};
  assign p2_sub_35099_comb = {p2_add_35033_comb, p2_umul_34248_comb[1:0]} - {p2_add_35035_comb, p2_umul_34063_comb[1:0]};
  assign p2_add_34242_comb = p2_umul_34112_comb[31:3] + p2_umul_34113_comb[31:3];
  assign p2_add_34244_comb = p2_umul_34197_comb + p2_concat_34198_comb;
  assign p2_add_34245_comb = p2_umul_34199_comb + p2_umul_34021_comb;
  assign p2_add_34306_comb = p2_umul_34200_comb[31:3] + p2_umul_34201_comb[31:3];
  assign p2_add_34308_comb = p2_umul_34248_comb + p2_concat_34249_comb;
  assign p2_add_34309_comb = p2_umul_34250_comb + p2_umul_34063_comb;
  assign p2_add_34754_comb = p2_umul_34600_comb[31:2] + p2_add_34605_comb;
  assign p2_sub_34755_comb = p2_or_34692_comb - p2_umul_34693_comb;
  assign p2_sub_34756_comb = p2_or_34692_comb - p2_umul_34694_comb;
  assign p2_sub_34757_comb = {p2_add_34605_comb, p2_umul_34467_comb[1:0]} - p2_umul_34696_comb;
  assign p2_add_34766_comb = p2_umul_34624_comb[31:2] + p2_add_34629_comb;
  assign p2_sub_34767_comb = p2_or_34710_comb - p2_umul_34711_comb;
  assign p2_sub_34768_comb = p2_or_34710_comb - p2_umul_34712_comb;
  assign p2_sub_34769_comb = {p2_add_34629_comb, p2_umul_34476_comb[1:0]} - p2_umul_34714_comb;
  assign p2_add_34770_comb = p2_umul_34632_comb[31:2] + p2_add_34637_comb;
  assign p2_sub_34771_comb = p2_or_34716_comb - p2_umul_34717_comb;
  assign p2_sub_34772_comb = p2_or_34716_comb - p2_umul_34718_comb;
  assign p2_sub_34773_comb = {p2_add_34637_comb, p2_umul_34479_comb[1:0]} - p2_umul_34720_comb;
  assign p2_add_34782_comb = p2_umul_34656_comb[31:2] + p2_add_34661_comb;
  assign p2_sub_34783_comb = p2_or_34734_comb - p2_umul_34735_comb;
  assign p2_sub_34784_comb = p2_or_34734_comb - p2_umul_34736_comb;
  assign p2_sub_34785_comb = {p2_add_34661_comb, p2_umul_34488_comb[1:0]} - p2_umul_34738_comb;
  assign p2_bit_slice_34411_comb = p2_sub_34349_comb[31:8];
  assign p2_bit_slice_34412_comb = p2_sub_34350_comb[31:8];
  assign p2_add_34413_comb = p2_sign_ext_34351_comb + p2_sign_ext_34352_comb;
  assign p2_bit_slice_34415_comb = p2_sub_34353_comb[31:8];
  assign p2_bit_slice_34416_comb = p2_sub_34354_comb[31:8];
  assign p2_add_34417_comb = p2_sign_ext_34355_comb + p2_sign_ext_34356_comb;
  assign p2_bit_slice_34423_comb = p2_sub_34361_comb[31:8];
  assign p2_bit_slice_34424_comb = p2_sub_34362_comb[31:8];
  assign p2_add_34425_comb = p2_sign_ext_34363_comb + p2_sign_ext_34364_comb;
  assign p2_bit_slice_34427_comb = p2_sub_34365_comb[31:8];
  assign p2_bit_slice_34428_comb = p2_sub_34366_comb[31:8];
  assign p2_add_34429_comb = p2_sign_ext_34367_comb + p2_sign_ext_34368_comb;
  assign p2_concat_35127_comb = {p2_add_35108_comb, p2_add_34997_comb[2:1]};
  assign p2_add_35114_comb = p2_sub_35064_comb[31:13] + 19'h0_0001;
  assign p2_bit_slice_35115_comb = p2_sub_35064_comb[12:8];
  assign p2_concat_35128_comb = {p2_add_35110_comb, p2_add_35002_comb[2:1]};
  assign p2_add_35117_comb = p2_sub_35067_comb[31:13] + 19'h0_0001;
  assign p2_bit_slice_35118_comb = p2_sub_35067_comb[12:8];
  assign p2_concat_35129_comb = {p2_add_35112_comb, p2_add_35007_comb[2:1]};
  assign p2_add_35120_comb = p2_sub_35070_comb[31:13] + 19'h0_0001;
  assign p2_bit_slice_35121_comb = p2_sub_35070_comb[12:8];
  assign p2_bit_slice_34799_comb = p2_add_34754_comb[29:1];
  assign p2_bit_slice_34800_comb = p2_sub_34755_comb[31:3];
  assign p2_bit_slice_34801_comb = p2_sub_34756_comb[31:3];
  assign p2_bit_slice_34802_comb = p2_sub_34757_comb[31:3];
  assign p2_bit_slice_34811_comb = p2_add_34766_comb[29:1];
  assign p2_bit_slice_34812_comb = p2_sub_34767_comb[31:3];
  assign p2_bit_slice_34813_comb = p2_sub_34768_comb[31:3];
  assign p2_bit_slice_34814_comb = p2_sub_34769_comb[31:3];
  assign p2_bit_slice_34815_comb = p2_add_34770_comb[29:1];
  assign p2_bit_slice_34816_comb = p2_sub_34771_comb[31:3];
  assign p2_bit_slice_34817_comb = p2_sub_34772_comb[31:3];
  assign p2_bit_slice_34818_comb = p2_sub_34773_comb[31:3];
  assign p2_bit_slice_34827_comb = p2_add_34782_comb[29:1];
  assign p2_bit_slice_34828_comb = p2_sub_34783_comb[31:3];
  assign p2_bit_slice_34829_comb = p2_sub_34784_comb[31:3];
  assign p2_bit_slice_34830_comb = p2_sub_34785_comb[31:3];
  assign p2_sign_ext_34468_comb = {{8{p2_bit_slice_34411_comb[23]}}, p2_bit_slice_34411_comb};
  assign p2_sign_ext_34469_comb = {{8{p2_bit_slice_34412_comb[23]}}, p2_bit_slice_34412_comb};
  assign p2_umul_34470_comb = umul32b_32b_x_10b(p2_add_34413_comb, 10'h235);
  assign p2_sign_ext_34471_comb = {{8{p2_bit_slice_34415_comb[23]}}, p2_bit_slice_34415_comb};
  assign p2_sign_ext_34472_comb = {{8{p2_bit_slice_34416_comb[23]}}, p2_bit_slice_34416_comb};
  assign p2_umul_34473_comb = umul32b_32b_x_10b(p2_add_34417_comb, 10'h235);
  assign p2_sign_ext_34480_comb = {{8{p2_bit_slice_34423_comb[23]}}, p2_bit_slice_34423_comb};
  assign p2_sign_ext_34481_comb = {{8{p2_bit_slice_34424_comb[23]}}, p2_bit_slice_34424_comb};
  assign p2_umul_34482_comb = umul32b_32b_x_10b(p2_add_34425_comb, 10'h235);
  assign p2_sign_ext_34483_comb = {{8{p2_bit_slice_34427_comb[23]}}, p2_bit_slice_34427_comb};
  assign p2_sign_ext_34484_comb = {{8{p2_bit_slice_34428_comb[23]}}, p2_bit_slice_34428_comb};
  assign p2_umul_34485_comb = umul32b_32b_x_10b(p2_add_34429_comb, 10'h235);
  assign p2_add_34433_comb = p2_sign_ext_34334_comb[31:7] + 25'h000_0001;
  assign p2_add_34435_comb = p1_umul_33520[31:11] + p1_bit_slice_33594;
  assign p2_add_34437_comb = p2_sign_ext_34335_comb[31:7] + 25'h000_0001;
  assign p2_add_34439_comb = p1_umul_33522[31:11] + p1_bit_slice_33596;
  assign p2_add_34441_comb = p2_sign_ext_34336_comb[31:7] + 25'h000_0001;
  assign p2_add_34443_comb = p1_umul_33591[31:11] + p1_bit_slice_33594;
  assign p2_add_34445_comb = p2_sign_ext_34337_comb[31:7] + 25'h000_0001;
  assign p2_add_34447_comb = p1_umul_33592[31:11] + p1_bit_slice_33596;
  assign p2_add_34449_comb = p1_umul_33591[31:7] + 25'h000_0001;
  assign p2_add_34450_comb = p2_sign_ext_34336_comb[31:2] + p1_umul_33520[31:2];
  assign p2_add_34451_comb = p1_umul_33592[31:7] + 25'h000_0001;
  assign p2_add_34452_comb = p2_sign_ext_34337_comb[31:2] + p1_umul_33522[31:2];
  assign p2_add_34453_comb = p1_umul_33520[31:7] + 25'h000_0001;
  assign p2_add_34454_comb = p2_sign_ext_34334_comb[31:3] + p1_umul_33591[31:3];
  assign p2_add_34455_comb = p1_umul_33522[31:7] + 25'h000_0001;
  assign p2_add_34456_comb = p2_sign_ext_34335_comb[31:3] + p1_umul_33592[31:3];
  assign p2_sign_ext_35136_comb = {{3{p2_concat_35127_comb[28]}}, p2_concat_35127_comb};
  assign p2_bit_slice_35116_comb = p2_sub_35093_comb[31:8];
  assign p2_sign_ext_35138_comb = {{3{p2_concat_35128_comb[28]}}, p2_concat_35128_comb};
  assign p2_bit_slice_35119_comb = p2_sub_35096_comb[31:8];
  assign p2_sign_ext_35140_comb = {{3{p2_concat_35129_comb[28]}}, p2_concat_35129_comb};
  assign p2_bit_slice_35122_comb = p2_sub_35099_comb[31:8];
  assign p2_add_35142_comb = p2_sub_35093_comb[31:13] + 19'h0_0001;
  assign p2_add_35144_comb = p2_sub_35096_comb[31:13] + 19'h0_0001;
  assign p2_add_35146_comb = p2_sub_35099_comb[31:13] + 19'h0_0001;
  assign p2_add_34338_comb = p2_add_34242_comb + p2_umul_34112_comb[31:3];
  assign p2_add_34340_comb = {p2_add_34242_comb, p2_umul_34113_comb[2:1]} + p2_add_34244_comb[31:1];
  assign p2_add_34342_comb = p2_add_34245_comb[31:3] + p2_umul_34112_comb[31:3];
  assign p2_add_34401_comb = p2_add_34306_comb + p2_umul_34200_comb[31:3];
  assign p2_add_34405_comb = {p2_add_34306_comb, p2_umul_34201_comb[2:1]} + p2_add_34308_comb[31:1];
  assign p2_add_34407_comb = p2_add_34309_comb[31:3] + p2_umul_34200_comb[31:3];
  assign p2_sign_ext_34853_comb = {{3{p2_bit_slice_34799_comb[28]}}, p2_bit_slice_34799_comb};
  assign p2_sign_ext_34854_comb = {{3{p2_bit_slice_34800_comb[28]}}, p2_bit_slice_34800_comb};
  assign p2_sign_ext_34855_comb = {{3{p2_bit_slice_34801_comb[28]}}, p2_bit_slice_34801_comb};
  assign p2_sign_ext_34856_comb = {{3{p2_bit_slice_34802_comb[28]}}, p2_bit_slice_34802_comb};
  assign p2_sign_ext_34857_comb = {{3{p2_bit_slice_34811_comb[28]}}, p2_bit_slice_34811_comb};
  assign p2_sign_ext_34858_comb = {{3{p2_bit_slice_34812_comb[28]}}, p2_bit_slice_34812_comb};
  assign p2_sign_ext_34859_comb = {{3{p2_bit_slice_34813_comb[28]}}, p2_bit_slice_34813_comb};
  assign p2_sign_ext_34860_comb = {{3{p2_bit_slice_34814_comb[28]}}, p2_bit_slice_34814_comb};
  assign p2_sign_ext_34861_comb = {{3{p2_bit_slice_34815_comb[28]}}, p2_bit_slice_34815_comb};
  assign p2_sign_ext_34862_comb = {{3{p2_bit_slice_34816_comb[28]}}, p2_bit_slice_34816_comb};
  assign p2_sign_ext_34863_comb = {{3{p2_bit_slice_34817_comb[28]}}, p2_bit_slice_34817_comb};
  assign p2_sign_ext_34864_comb = {{3{p2_bit_slice_34818_comb[28]}}, p2_bit_slice_34818_comb};
  assign p2_sign_ext_34865_comb = {{3{p2_bit_slice_34827_comb[28]}}, p2_bit_slice_34827_comb};
  assign p2_sign_ext_34866_comb = {{3{p2_bit_slice_34828_comb[28]}}, p2_bit_slice_34828_comb};
  assign p2_sign_ext_34867_comb = {{3{p2_bit_slice_34829_comb[28]}}, p2_bit_slice_34829_comb};
  assign p2_sign_ext_34868_comb = {{3{p2_bit_slice_34830_comb[28]}}, p2_bit_slice_34830_comb};
  assign p2_add_34517_comb = p2_sign_ext_34468_comb + p2_sign_ext_34469_comb;
  assign p2_add_34522_comb = p2_sign_ext_34471_comb + p2_sign_ext_34472_comb;
  assign p2_add_34537_comb = p2_sign_ext_34480_comb + p2_sign_ext_34481_comb;
  assign p2_add_34542_comb = p2_sign_ext_34483_comb + p2_sign_ext_34484_comb;
  assign p2_add_35149_comb = p2_bit_slice_35116_comb + {p2_add_35114_comb, p2_bit_slice_35115_comb};
  assign p2_add_35151_comb = p2_bit_slice_35119_comb + {p2_add_35117_comb, p2_bit_slice_35118_comb};
  assign p2_add_35153_comb = p2_bit_slice_35122_comb + {p2_add_35120_comb, p2_bit_slice_35121_comb};
  assign p2_bit_slice_35154_comb = p2_sub_35064_comb[31:8];
  assign p2_bit_slice_35155_comb = p2_sub_35067_comb[31:8];
  assign p2_bit_slice_35156_comb = p2_sub_35070_comb[31:8];
  assign p2_add_34399_comb = p2_add_34244_comb + p2_add_34245_comb;
  assign p2_add_34459_comb = p2_add_34308_comb + p2_add_34309_comb;
  assign p2_add_34908_comb = p2_sign_ext_34853_comb + p2_sign_ext_34854_comb;
  assign p2_add_34909_comb = p2_sign_ext_34855_comb + p2_sign_ext_34856_comb;
  assign p2_add_34910_comb = p2_sign_ext_34857_comb + p2_sign_ext_34858_comb;
  assign p2_add_34911_comb = p2_sign_ext_34859_comb + p2_sign_ext_34860_comb;
  assign p2_add_34912_comb = p2_sign_ext_34861_comb + p2_sign_ext_34862_comb;
  assign p2_add_34913_comb = p2_sign_ext_34863_comb + p2_sign_ext_34864_comb;
  assign p2_add_34914_comb = p2_sign_ext_34865_comb + p2_sign_ext_34866_comb;
  assign p2_add_34915_comb = p2_sign_ext_34867_comb + p2_sign_ext_34868_comb;
  assign p2_add_34995_comb = p2_sign_ext_34853_comb + p2_sign_ext_34856_comb;
  assign p2_add_34996_comb = p2_sign_ext_34855_comb + p2_sign_ext_34854_comb;
  assign p2_add_35000_comb = p2_sign_ext_34857_comb + p2_sign_ext_34860_comb;
  assign p2_add_35001_comb = p2_sign_ext_34859_comb + p2_sign_ext_34858_comb;
  assign p2_add_35005_comb = p2_sign_ext_34861_comb + p2_sign_ext_34864_comb;
  assign p2_add_35006_comb = p2_sign_ext_34863_comb + p2_sign_ext_34862_comb;
  assign p2_add_35010_comb = p2_sign_ext_34865_comb + p2_sign_ext_34868_comb;
  assign p2_add_35011_comb = p2_sign_ext_34867_comb + p2_sign_ext_34866_comb;
  assign p2_umul_34608_comb = umul32b_32b_x_12b(p2_sign_ext_34351_comb, 12'h8e4);
  assign p2_umul_34609_comb = umul32b_32b_x_12b(p2_add_34517_comb, 12'h968);
  assign p2_add_34613_comb = p2_umul_34470_comb[31:2] + 30'h0000_0001;
  assign p2_umul_34616_comb = umul32b_32b_x_12b(p2_sign_ext_34355_comb, 12'h8e4);
  assign p2_umul_34617_comb = umul32b_32b_x_12b(p2_add_34522_comb, 12'h968);
  assign p2_add_34621_comb = p2_umul_34473_comb[31:2] + 30'h0000_0001;
  assign p2_umul_34640_comb = umul32b_32b_x_12b(p2_sign_ext_34363_comb, 12'h8e4);
  assign p2_umul_34641_comb = umul32b_32b_x_12b(p2_add_34537_comb, 12'h968);
  assign p2_add_34645_comb = p2_umul_34482_comb[31:2] + 30'h0000_0001;
  assign p2_umul_34648_comb = umul32b_32b_x_12b(p2_sign_ext_34367_comb, 12'h8e4);
  assign p2_umul_34649_comb = umul32b_32b_x_12b(p2_add_34542_comb, 12'h968);
  assign p2_add_34653_comb = p2_umul_34485_comb[31:2] + 30'h0000_0001;
  assign p2_add_34551_comb = {p2_add_34433_comb, p2_add_34238_comb[7:3]} + {p2_add_34435_comb, p1_umul_33520[10:2]};
  assign p2_add_34553_comb = p1_umul_33591[31:11] + p1_bit_slice_33593;
  assign p2_add_34555_comb = {p2_add_34437_comb, p2_add_34239_comb[7:3]} + {p2_add_34439_comb, p1_umul_33522[10:2]};
  assign p2_add_34557_comb = p1_umul_33592[31:11] + p1_bit_slice_33595;
  assign p2_add_34559_comb = {p2_add_34441_comb, p2_add_34240_comb[7:4]} + {p2_add_34443_comb, p1_umul_33591[10:3]};
  assign p2_add_34561_comb = p1_umul_33520[31:11] + p1_bit_slice_33593;
  assign p2_add_34563_comb = {p2_add_34445_comb, p2_add_34241_comb[7:4]} + {p2_add_34447_comb, p1_umul_33592[10:3]};
  assign p2_add_34565_comb = p1_umul_33522[31:11] + p1_bit_slice_33595;
  assign p2_add_34567_comb = p2_add_34449_comb[24:4] + p1_bit_slice_33594;
  assign p2_add_34570_comb = p2_add_34450_comb[29:9] + p1_bit_slice_33593;
  assign p2_add_34573_comb = p2_add_34451_comb[24:4] + p1_bit_slice_33596;
  assign p2_add_34576_comb = p2_add_34452_comb[29:9] + p1_bit_slice_33595;
  assign p2_add_34579_comb = p2_add_34453_comb[24:4] + p1_bit_slice_33594;
  assign p2_add_34582_comb = p2_add_34454_comb[28:8] + p1_bit_slice_33593;
  assign p2_add_34585_comb = p2_add_34455_comb[24:4] + p1_bit_slice_33596;
  assign p2_add_34588_comb = p2_add_34456_comb[28:8] + p1_bit_slice_33595;
  assign p2_sub_34919_comb = p2_umul_34112_comb - p2_umul_34197_comb;
  assign p2_sub_34968_comb = p2_umul_34200_comb - p2_umul_34248_comb;
  assign p2_add_35163_comb = p2_sign_ext_35136_comb[31:8] + p2_add_35149_comb;
  assign p2_add_35165_comb = p2_sign_ext_35138_comb[31:8] + p2_add_35151_comb;
  assign p2_add_35167_comb = p2_sign_ext_35140_comb[31:8] + p2_add_35153_comb;
  assign p2_add_35173_comb = {p2_add_35142_comb, p2_sub_35093_comb[12:8]} + p2_bit_slice_35154_comb;
  assign p2_add_35175_comb = p2_sign_ext_34858_comb + p2_sign_ext_34860_comb;
  assign p2_add_35176_comb = {p2_add_35144_comb, p2_sub_35096_comb[12:8]} + p2_bit_slice_35155_comb;
  assign p2_add_35178_comb = p2_sign_ext_34862_comb + p2_sign_ext_34864_comb;
  assign p2_add_35179_comb = {p2_add_35146_comb, p2_sub_35099_comb[12:8]} + p2_bit_slice_35156_comb;
  assign p2_add_35181_comb = p2_sign_ext_34866_comb + p2_sign_ext_34868_comb;
  assign p2_sub_34457_comb = p2_add_34399_comb - {p2_add_34338_comb, p2_umul_34113_comb[2:0]};
  assign p2_sub_34461_comb = {p2_add_34340_comb, p2_add_34244_comb[0]} - {p2_add_34342_comb, p2_add_34245_comb[2:0]};
  assign p2_sub_34506_comb = p2_add_34459_comb - {p2_add_34401_comb, p2_umul_34201_comb[2:0]};
  assign p2_sub_34509_comb = {p2_add_34405_comb, p2_add_34308_comb[0]} - {p2_add_34407_comb, p2_add_34309_comb[2:0]};
  assign p2_sub_34951_comb = p2_add_34908_comb - p2_add_34909_comb;
  assign p2_sub_34953_comb = p2_add_34910_comb - p2_add_34911_comb;
  assign p2_sub_34955_comb = p2_add_34912_comb - p2_add_34913_comb;
  assign p2_sub_34957_comb = p2_add_34914_comb - p2_add_34915_comb;
  assign p2_sub_35044_comb = p2_add_34995_comb - p2_add_34996_comb;
  assign p2_sub_35048_comb = p2_add_35000_comb - p2_add_35001_comb;
  assign p2_sub_35052_comb = p2_add_35005_comb - p2_add_35006_comb;
  assign p2_sub_35056_comb = p2_add_35010_comb - p2_add_35011_comb;
  assign p2_or_34698_comb = p2_umul_34609_comb | 32'h0000_0004;
  assign p2_umul_34699_comb = umul32b_32b_x_12b(p2_sign_ext_34469_comb, 12'hfb1);
  assign p2_umul_34700_comb = umul32b_32b_x_10b(p2_sign_ext_34468_comb, 10'h31f);
  assign p2_umul_34702_comb = umul32b_32b_x_12b(p2_sign_ext_34352_comb, 12'hd4e);
  assign p2_or_34704_comb = p2_umul_34617_comb | 32'h0000_0004;
  assign p2_umul_34705_comb = umul32b_32b_x_12b(p2_sign_ext_34472_comb, 12'hfb1);
  assign p2_umul_34706_comb = umul32b_32b_x_10b(p2_sign_ext_34471_comb, 10'h31f);
  assign p2_umul_34708_comb = umul32b_32b_x_12b(p2_sign_ext_34356_comb, 12'hd4e);
  assign p2_or_34722_comb = p2_umul_34641_comb | 32'h0000_0004;
  assign p2_umul_34723_comb = umul32b_32b_x_12b(p2_sign_ext_34481_comb, 12'hfb1);
  assign p2_umul_34724_comb = umul32b_32b_x_10b(p2_sign_ext_34480_comb, 10'h31f);
  assign p2_umul_34726_comb = umul32b_32b_x_12b(p2_sign_ext_34364_comb, 12'hd4e);
  assign p2_or_34728_comb = p2_umul_34649_comb | 32'h0000_0004;
  assign p2_umul_34729_comb = umul32b_32b_x_12b(p2_sign_ext_34484_comb, 12'hfb1);
  assign p2_umul_34730_comb = umul32b_32b_x_10b(p2_sign_ext_34483_comb, 10'h31f);
  assign p2_umul_34732_comb = umul32b_32b_x_12b(p2_sign_ext_34368_comb, 12'hd4e);
  assign p2_add_34965_comb = p2_sub_34919_comb + p2_concat_34198_comb;
  assign p2_add_34966_comb = p2_add_34796_comb[26:2] + {p2_add_34841_comb, 4'h1};
  assign p2_add_35017_comb = p2_sub_34968_comb + p2_concat_34249_comb;
  assign p2_add_35018_comb = p2_add_34852_comb[26:2] + {p2_add_34885_comb, 4'h1};
  assign p2_add_35183_comb = p2_sign_ext_34859_comb + p2_sign_ext_34857_comb;
  assign p2_concat_35184_comb = {p2_add_35163_comb, p2_add_35108_comb[5:0], p2_add_34997_comb[2:1]};
  assign p2_add_35185_comb = p2_sign_ext_34863_comb + p2_sign_ext_34861_comb;
  assign p2_concat_35186_comb = {p2_add_35165_comb, p2_add_35110_comb[5:0], p2_add_35002_comb[2:1]};
  assign p2_add_35187_comb = p2_sign_ext_34867_comb + p2_sign_ext_34865_comb;
  assign p2_concat_35188_comb = {p2_add_35167_comb, p2_add_35112_comb[5:0], p2_add_35007_comb[2:1]};
  assign p2_sub_35189_comb = {p2_add_35149_comb, 8'h00} - p2_sign_ext_35136_comb;
  assign p2_sub_35190_comb = {p2_add_35151_comb, 8'h00} - p2_sign_ext_35138_comb;
  assign p2_sub_35191_comb = {p2_add_35153_comb, 8'h00} - p2_sign_ext_35140_comb;
  assign p2_add_35193_comb = p2_sign_ext_35136_comb + p2_add_35175_comb;
  assign p2_add_35195_comb = p2_sign_ext_35138_comb + p2_add_35178_comb;
  assign p2_add_35197_comb = p2_sign_ext_35140_comb + p2_add_35181_comb;
  assign p2_umul_34505_comb = umul32b_32b_x_8b(p2_sub_34457_comb, 8'hb5);
  assign p2_umul_34508_comb = umul32b_32b_x_8b(p2_sub_34461_comb, 8'hb5);
  assign p2_umul_34593_comb = umul32b_32b_x_8b(p2_sub_34506_comb, 8'hb5);
  assign p2_umul_34596_comb = umul32b_32b_x_8b(p2_sub_34509_comb, 8'hb5);
  assign p2_umul_34991_comb = umul32b_32b_x_8b(p2_sub_34951_comb, 8'hb5);
  assign p2_umul_34992_comb = umul32b_32b_x_8b(p2_sub_34953_comb, 8'hb5);
  assign p2_umul_34993_comb = umul32b_32b_x_8b(p2_sub_34955_comb, 8'hb5);
  assign p2_umul_34994_comb = umul32b_32b_x_8b(p2_sub_34957_comb, 8'hb5);
  assign p2_umul_35077_comb = umul32b_32b_x_8b(p2_sub_35044_comb, 8'hb5);
  assign p2_umul_35079_comb = umul32b_32b_x_8b(p2_sub_35048_comb, 8'hb5);
  assign p2_umul_35081_comb = umul32b_32b_x_8b(p2_sub_35052_comb, 8'hb5);
  assign p2_umul_35083_comb = umul32b_32b_x_8b(p2_sub_35056_comb, 8'hb5);
  assign p2_add_34758_comb = p2_umul_34608_comb[31:2] + p2_add_34613_comb;
  assign p2_sub_34759_comb = p2_or_34698_comb - p2_umul_34699_comb;
  assign p2_sub_34760_comb = p2_or_34698_comb - p2_umul_34700_comb;
  assign p2_sub_34761_comb = {p2_add_34613_comb, p2_umul_34470_comb[1:0]} - p2_umul_34702_comb;
  assign p2_add_34762_comb = p2_umul_34616_comb[31:2] + p2_add_34621_comb;
  assign p2_sub_34763_comb = p2_or_34704_comb - p2_umul_34705_comb;
  assign p2_sub_34764_comb = p2_or_34704_comb - p2_umul_34706_comb;
  assign p2_sub_34765_comb = {p2_add_34621_comb, p2_umul_34473_comb[1:0]} - p2_umul_34708_comb;
  assign p2_add_34774_comb = p2_umul_34640_comb[31:2] + p2_add_34645_comb;
  assign p2_sub_34775_comb = p2_or_34722_comb - p2_umul_34723_comb;
  assign p2_sub_34776_comb = p2_or_34722_comb - p2_umul_34724_comb;
  assign p2_sub_34777_comb = {p2_add_34645_comb, p2_umul_34482_comb[1:0]} - p2_umul_34726_comb;
  assign p2_add_34778_comb = p2_umul_34648_comb[31:2] + p2_add_34653_comb;
  assign p2_sub_34779_comb = p2_or_34728_comb - p2_umul_34729_comb;
  assign p2_sub_34780_comb = p2_or_34728_comb - p2_umul_34730_comb;
  assign p2_sub_34781_comb = {p2_add_34653_comb, p2_umul_34485_comb[1:0]} - p2_umul_34732_comb;
  assign p2_sub_34739_comb = {p2_add_34551_comb, p2_add_34238_comb[2:1]} - {p2_add_34553_comb, p1_umul_33591[10:0]};
  assign p2_sub_34740_comb = {p2_add_34555_comb, p2_add_34239_comb[2:1]} - {p2_add_34557_comb, p1_umul_33592[10:0]};
  assign p2_sub_34741_comb = {p2_add_34559_comb, p2_add_34240_comb[3:1]} - {p2_add_34561_comb, p1_umul_33520[10:0]};
  assign p2_sub_34742_comb = {p2_add_34563_comb, p2_add_34241_comb[3:1]} - {p2_add_34565_comb, p1_umul_33522[10:0]};
  assign p2_sub_34743_comb = {p2_add_34567_comb, p2_add_34449_comb[3:0], p1_umul_33591[6:0]} - {p2_add_34570_comb, p2_add_34450_comb[8:0], p2_add_34240_comb[2:1]};
  assign p2_sub_34744_comb = {p2_add_34573_comb, p2_add_34451_comb[3:0], p1_umul_33592[6:0]} - {p2_add_34576_comb, p2_add_34452_comb[8:0], p2_add_34241_comb[2:1]};
  assign p2_sub_34745_comb = {p2_add_34579_comb, p2_add_34453_comb[3:0], p1_umul_33520[6:0]} - {p2_add_34582_comb, p2_add_34454_comb[7:0], p2_add_34238_comb[3:1]};
  assign p2_sub_34746_comb = {p2_add_34585_comb, p2_add_34455_comb[3:0], p1_umul_33522[6:0]} - {p2_add_34588_comb, p2_add_34456_comb[7:0], p2_add_34239_comb[3:1]};
  assign p2_umul_35047_comb = umul32b_32b_x_12b(p2_sign_ext_34832_comb, 12'hec8);
  assign p2_umul_35051_comb = umul32b_32b_x_12b(p2_sign_ext_34834_comb, 12'hec8);
  assign p2_umul_35055_comb = umul32b_32b_x_12b(p2_sign_ext_34836_comb, 12'hec8);
  assign p2_add_35198_comb = p2_add_35183_comb + p2_concat_35184_comb;
  assign p2_add_35199_comb = p2_add_35185_comb + p2_concat_35186_comb;
  assign p2_add_35200_comb = p2_add_35187_comb + p2_concat_35188_comb;
  assign p2_add_35201_comb = p2_sub_35189_comb + p2_add_35175_comb;
  assign p2_add_35202_comb = p2_sub_35190_comb + p2_add_35178_comb;
  assign p2_add_35203_comb = p2_sub_35191_comb + p2_add_35181_comb;
  assign p2_sub_35204_comb = {p2_add_35173_comb, 8'h00} - p2_add_35193_comb;
  assign p2_sub_35205_comb = {p2_add_35176_comb, 8'h00} - p2_add_35195_comb;
  assign p2_sub_35206_comb = {p2_add_35179_comb, 8'h00} - p2_add_35197_comb;
  assign p2_sub_35207_comb = p2_concat_35184_comb - p2_add_35183_comb;
  assign p2_sub_35208_comb = p2_concat_35186_comb - p2_add_35185_comb;
  assign p2_sub_35209_comb = p2_concat_35188_comb - p2_add_35187_comb;
  assign p2_bit_slice_34803_comb = p2_add_34758_comb[29:1];
  assign p2_bit_slice_34804_comb = p2_sub_34759_comb[31:3];
  assign p2_bit_slice_34805_comb = p2_sub_34760_comb[31:3];
  assign p2_bit_slice_34806_comb = p2_sub_34761_comb[31:3];
  assign p2_bit_slice_34807_comb = p2_add_34762_comb[29:1];
  assign p2_bit_slice_34808_comb = p2_sub_34763_comb[31:3];
  assign p2_bit_slice_34809_comb = p2_sub_34764_comb[31:3];
  assign p2_bit_slice_34810_comb = p2_sub_34765_comb[31:3];
  assign p2_bit_slice_34819_comb = p2_add_34774_comb[29:1];
  assign p2_bit_slice_34820_comb = p2_sub_34775_comb[31:3];
  assign p2_bit_slice_34821_comb = p2_sub_34776_comb[31:3];
  assign p2_bit_slice_34822_comb = p2_sub_34777_comb[31:3];
  assign p2_bit_slice_34823_comb = p2_add_34778_comb[29:1];
  assign p2_bit_slice_34824_comb = p2_sub_34779_comb[31:3];
  assign p2_bit_slice_34825_comb = p2_sub_34780_comb[31:3];
  assign p2_bit_slice_34826_comb = p2_sub_34781_comb[31:3];
  assign p2_bit_slice_34786_comb = p2_sub_34739_comb[31:8];
  assign p2_bit_slice_34787_comb = p2_sub_34740_comb[31:8];
  assign p2_bit_slice_34788_comb = p2_sub_34741_comb[31:8];
  assign p2_bit_slice_34789_comb = p2_sub_34742_comb[31:8];
  assign p2_bit_slice_34790_comb = p2_sub_34743_comb[31:8];
  assign p2_bit_slice_34791_comb = p2_sub_34744_comb[31:8];
  assign p2_bit_slice_34792_comb = p2_sub_34745_comb[31:8];
  assign p2_bit_slice_34793_comb = p2_sub_34746_comb[31:8];
  assign p2_add_35061_comb = p2_add_34965_comb[31:2] + {p2_add_34966_comb, p2_add_34796_comb[1:0], p2_umul_34687_comb[4:2]};
  assign p2_sub_35078_comb = {p2_add_34997_comb, 2'h0} - p2_umul_35047_comb;
  assign p2_sub_35080_comb = {p2_add_35002_comb, 2'h0} - p2_umul_35051_comb;
  assign p2_sub_35082_comb = {p2_add_35007_comb, 2'h0} - p2_umul_35055_comb;
  assign p2_add_35090_comb = p2_add_35017_comb[31:2] + {p2_add_35018_comb, p2_add_34852_comb[1:0], p2_umul_34753_comb[4:2]};
  assign p2_add_35172_comb = p2_sign_ext_34854_comb + p2_sign_ext_34856_comb;
  assign p2_add_35182_comb = p2_sign_ext_34855_comb + p2_sign_ext_34853_comb;
  assign p2_bit_slice_35210_comb = p2_add_35198_comb[31:14];
  assign p2_bit_slice_35211_comb = p2_add_35199_comb[31:14];
  assign p2_bit_slice_35212_comb = p2_add_35200_comb[31:14];
  assign p2_bit_slice_35213_comb = p2_add_35201_comb[31:14];
  assign p2_bit_slice_35214_comb = p2_add_35202_comb[31:14];
  assign p2_bit_slice_35215_comb = p2_add_35203_comb[31:14];
  assign p2_bit_slice_35216_comb = p2_sub_35204_comb[31:14];
  assign p2_bit_slice_35217_comb = p2_sub_35205_comb[31:14];
  assign p2_bit_slice_35218_comb = p2_sub_35206_comb[31:14];
  assign p2_bit_slice_35219_comb = p2_sub_35207_comb[31:14];
  assign p2_bit_slice_35220_comb = p2_sub_35208_comb[31:14];
  assign p2_bit_slice_35221_comb = p2_sub_35209_comb[31:14];
  assign p2_add_34680_comb = p2_umul_34505_comb[31:7] + 25'h000_0001;
  assign p2_add_34683_comb = p2_umul_34508_comb[31:7] + 25'h000_0001;
  assign p2_add_34747_comb = p2_umul_34593_comb[31:7] + 25'h000_0001;
  assign p2_add_34749_comb = p2_umul_34596_comb[31:7] + 25'h000_0001;
  assign p2_add_35073_comb = p2_umul_34991_comb[31:7] + 25'h000_0001;
  assign p2_add_35074_comb = p2_umul_34992_comb[31:7] + 25'h000_0001;
  assign p2_add_35075_comb = p2_umul_34993_comb[31:7] + 25'h000_0001;
  assign p2_add_35076_comb = p2_umul_34994_comb[31:7] + 25'h000_0001;
  assign p2_add_35123_comb = p2_umul_35077_comb[31:7] + 25'h000_0001;
  assign p2_add_35124_comb = p2_umul_35079_comb[31:7] + 25'h000_0001;
  assign p2_add_35125_comb = p2_umul_35081_comb[31:7] + 25'h000_0001;
  assign p2_add_35126_comb = p2_umul_35083_comb[31:7] + 25'h000_0001;
  assign p2_umul_34794_comb = umul32b_32b_x_12b(p1_array_index_33710, 12'hec8);
  assign p2_umul_34837_comb = umul32b_32b_x_12b(p1_array_index_33740, 12'hec8);

  // Registers for pipe stage 2:
  reg [28:0] p2_bit_slice_34803;
  reg [28:0] p2_bit_slice_34804;
  reg [28:0] p2_bit_slice_34805;
  reg [28:0] p2_bit_slice_34806;
  reg [28:0] p2_bit_slice_34807;
  reg [28:0] p2_bit_slice_34808;
  reg [28:0] p2_bit_slice_34809;
  reg [28:0] p2_bit_slice_34810;
  reg [28:0] p2_bit_slice_34819;
  reg [28:0] p2_bit_slice_34820;
  reg [28:0] p2_bit_slice_34821;
  reg [28:0] p2_bit_slice_34822;
  reg [28:0] p2_bit_slice_34823;
  reg [28:0] p2_bit_slice_34824;
  reg [28:0] p2_bit_slice_34825;
  reg [28:0] p2_bit_slice_34826;
  reg [23:0] p2_bit_slice_33771;
  reg [23:0] p2_bit_slice_33772;
  reg [23:0] p2_bit_slice_34786;
  reg [23:0] p2_bit_slice_34787;
  reg [23:0] p2_bit_slice_34788;
  reg [23:0] p2_bit_slice_34789;
  reg [23:0] p2_bit_slice_34790;
  reg [23:0] p2_bit_slice_34791;
  reg [23:0] p2_bit_slice_34792;
  reg [23:0] p2_bit_slice_34793;
  reg [20:0] p2_bit_slice_33779;
  reg [20:0] p2_bit_slice_33780;
  reg [20:0] p2_bit_slice_33783;
  reg [20:0] p2_bit_slice_33784;
  reg [29:0] p2_add_35061;
  reg [31:0] p2_sub_35078;
  reg [31:0] p2_sub_35080;
  reg [31:0] p2_sub_35082;
  reg [29:0] p2_add_35090;
  reg [4:0] p2_bit_slice_35115;
  reg [23:0] p2_bit_slice_35116;
  reg [4:0] p2_bit_slice_35118;
  reg [23:0] p2_bit_slice_35119;
  reg [4:0] p2_bit_slice_35121;
  reg [23:0] p2_bit_slice_35122;
  reg [23:0] p2_bit_slice_35154;
  reg [23:0] p2_bit_slice_35155;
  reg [23:0] p2_bit_slice_35156;
  reg [31:0] p2_add_35172;
  reg [31:0] p2_add_35182;
  reg [17:0] p2_bit_slice_35210;
  reg [17:0] p2_bit_slice_35211;
  reg [17:0] p2_bit_slice_35212;
  reg [17:0] p2_bit_slice_35213;
  reg [17:0] p2_bit_slice_35214;
  reg [17:0] p2_bit_slice_35215;
  reg [17:0] p2_bit_slice_35216;
  reg [17:0] p2_bit_slice_35217;
  reg [17:0] p2_bit_slice_35218;
  reg [17:0] p2_bit_slice_35219;
  reg [17:0] p2_bit_slice_35220;
  reg [17:0] p2_bit_slice_35221;
  reg [24:0] p2_add_34680;
  reg [24:0] p2_add_34683;
  reg [24:0] p2_add_34747;
  reg [24:0] p2_add_34749;
  reg [24:0] p2_add_35073;
  reg [24:0] p2_add_35074;
  reg [24:0] p2_add_35075;
  reg [24:0] p2_add_35076;
  reg [18:0] p2_add_35114;
  reg [18:0] p2_add_35117;
  reg [18:0] p2_add_35120;
  reg [24:0] p2_add_35123;
  reg [24:0] p2_add_35124;
  reg [24:0] p2_add_35125;
  reg [24:0] p2_add_35126;
  reg [31:0] p2_umul_34687;
  reg [31:0] p2_umul_34753;
  reg [31:0] p2_umul_34794;
  reg [31:0] p2_umul_34837;
  always_ff @ (posedge clk) begin
    p2_bit_slice_34803 <= p2_bit_slice_34803_comb;
    p2_bit_slice_34804 <= p2_bit_slice_34804_comb;
    p2_bit_slice_34805 <= p2_bit_slice_34805_comb;
    p2_bit_slice_34806 <= p2_bit_slice_34806_comb;
    p2_bit_slice_34807 <= p2_bit_slice_34807_comb;
    p2_bit_slice_34808 <= p2_bit_slice_34808_comb;
    p2_bit_slice_34809 <= p2_bit_slice_34809_comb;
    p2_bit_slice_34810 <= p2_bit_slice_34810_comb;
    p2_bit_slice_34819 <= p2_bit_slice_34819_comb;
    p2_bit_slice_34820 <= p2_bit_slice_34820_comb;
    p2_bit_slice_34821 <= p2_bit_slice_34821_comb;
    p2_bit_slice_34822 <= p2_bit_slice_34822_comb;
    p2_bit_slice_34823 <= p2_bit_slice_34823_comb;
    p2_bit_slice_34824 <= p2_bit_slice_34824_comb;
    p2_bit_slice_34825 <= p2_bit_slice_34825_comb;
    p2_bit_slice_34826 <= p2_bit_slice_34826_comb;
    p2_bit_slice_33771 <= p1_bit_slice_33771;
    p2_bit_slice_33772 <= p1_bit_slice_33772;
    p2_bit_slice_34786 <= p2_bit_slice_34786_comb;
    p2_bit_slice_34787 <= p2_bit_slice_34787_comb;
    p2_bit_slice_34788 <= p2_bit_slice_34788_comb;
    p2_bit_slice_34789 <= p2_bit_slice_34789_comb;
    p2_bit_slice_34790 <= p2_bit_slice_34790_comb;
    p2_bit_slice_34791 <= p2_bit_slice_34791_comb;
    p2_bit_slice_34792 <= p2_bit_slice_34792_comb;
    p2_bit_slice_34793 <= p2_bit_slice_34793_comb;
    p2_bit_slice_33779 <= p1_bit_slice_33779;
    p2_bit_slice_33780 <= p1_bit_slice_33780;
    p2_bit_slice_33783 <= p1_bit_slice_33783;
    p2_bit_slice_33784 <= p1_bit_slice_33784;
    p2_add_35061 <= p2_add_35061_comb;
    p2_sub_35078 <= p2_sub_35078_comb;
    p2_sub_35080 <= p2_sub_35080_comb;
    p2_sub_35082 <= p2_sub_35082_comb;
    p2_add_35090 <= p2_add_35090_comb;
    p2_bit_slice_35115 <= p2_bit_slice_35115_comb;
    p2_bit_slice_35116 <= p2_bit_slice_35116_comb;
    p2_bit_slice_35118 <= p2_bit_slice_35118_comb;
    p2_bit_slice_35119 <= p2_bit_slice_35119_comb;
    p2_bit_slice_35121 <= p2_bit_slice_35121_comb;
    p2_bit_slice_35122 <= p2_bit_slice_35122_comb;
    p2_bit_slice_35154 <= p2_bit_slice_35154_comb;
    p2_bit_slice_35155 <= p2_bit_slice_35155_comb;
    p2_bit_slice_35156 <= p2_bit_slice_35156_comb;
    p2_add_35172 <= p2_add_35172_comb;
    p2_add_35182 <= p2_add_35182_comb;
    p2_bit_slice_35210 <= p2_bit_slice_35210_comb;
    p2_bit_slice_35211 <= p2_bit_slice_35211_comb;
    p2_bit_slice_35212 <= p2_bit_slice_35212_comb;
    p2_bit_slice_35213 <= p2_bit_slice_35213_comb;
    p2_bit_slice_35214 <= p2_bit_slice_35214_comb;
    p2_bit_slice_35215 <= p2_bit_slice_35215_comb;
    p2_bit_slice_35216 <= p2_bit_slice_35216_comb;
    p2_bit_slice_35217 <= p2_bit_slice_35217_comb;
    p2_bit_slice_35218 <= p2_bit_slice_35218_comb;
    p2_bit_slice_35219 <= p2_bit_slice_35219_comb;
    p2_bit_slice_35220 <= p2_bit_slice_35220_comb;
    p2_bit_slice_35221 <= p2_bit_slice_35221_comb;
    p2_add_34680 <= p2_add_34680_comb;
    p2_add_34683 <= p2_add_34683_comb;
    p2_add_34747 <= p2_add_34747_comb;
    p2_add_34749 <= p2_add_34749_comb;
    p2_add_35073 <= p2_add_35073_comb;
    p2_add_35074 <= p2_add_35074_comb;
    p2_add_35075 <= p2_add_35075_comb;
    p2_add_35076 <= p2_add_35076_comb;
    p2_add_35114 <= p2_add_35114_comb;
    p2_add_35117 <= p2_add_35117_comb;
    p2_add_35120 <= p2_add_35120_comb;
    p2_add_35123 <= p2_add_35123_comb;
    p2_add_35124 <= p2_add_35124_comb;
    p2_add_35125 <= p2_add_35125_comb;
    p2_add_35126 <= p2_add_35126_comb;
    p2_umul_34687 <= p2_umul_34687_comb;
    p2_umul_34753 <= p2_umul_34753_comb;
    p2_umul_34794 <= p2_umul_34794_comb;
    p2_umul_34837 <= p2_umul_34837_comb;
  end

  // ===== Pipe stage 3:
  wire [23:0] p3_bit_slice_35376_comb;
  wire [23:0] p3_bit_slice_35377_comb;
  wire [31:0] p3_sign_ext_35378_comb;
  wire [23:0] p3_bit_slice_35379_comb;
  wire [31:0] p3_sign_ext_35380_comb;
  wire [23:0] p3_bit_slice_35381_comb;
  wire [31:0] p3_sign_ext_35382_comb;
  wire [31:0] p3_sign_ext_35383_comb;
  wire [31:0] p3_sign_ext_35384_comb;
  wire [31:0] p3_sign_ext_35385_comb;
  wire [31:0] p3_sign_ext_35386_comb;
  wire [31:0] p3_sign_ext_35387_comb;
  wire [31:0] p3_sign_ext_35388_comb;
  wire [31:0] p3_sign_ext_35389_comb;
  wire [31:0] p3_sign_ext_35390_comb;
  wire [31:0] p3_sign_ext_35391_comb;
  wire [31:0] p3_sign_ext_35395_comb;
  wire [31:0] p3_sign_ext_35399_comb;
  wire [31:0] p3_sign_ext_35408_comb;
  wire [31:0] p3_sign_ext_35409_comb;
  wire [31:0] p3_sign_ext_35410_comb;
  wire [31:0] p3_sign_ext_35411_comb;
  wire [31:0] p3_sign_ext_35412_comb;
  wire [31:0] p3_sign_ext_35413_comb;
  wire [31:0] p3_sign_ext_35414_comb;
  wire [31:0] p3_sign_ext_35415_comb;
  wire [31:0] p3_sign_ext_35416_comb;
  wire [31:0] p3_sign_ext_35417_comb;
  wire [31:0] p3_sign_ext_35418_comb;
  wire [31:0] p3_sign_ext_35419_comb;
  wire [31:0] p3_sign_ext_35420_comb;
  wire [31:0] p3_sign_ext_35421_comb;
  wire [31:0] p3_sign_ext_35422_comb;
  wire [31:0] p3_sign_ext_35423_comb;
  wire [31:0] p3_add_35424_comb;
  wire [31:0] p3_add_35426_comb;
  wire [31:0] p3_add_35428_comb;
  wire [31:0] p3_add_35430_comb;
  wire [31:0] p3_add_35432_comb;
  wire [24:0] p3_add_35434_comb;
  wire [20:0] p3_add_35436_comb;
  wire [24:0] p3_add_35441_comb;
  wire [20:0] p3_add_35443_comb;
  wire [24:0] p3_add_35448_comb;
  wire [29:0] p3_add_35449_comb;
  wire [24:0] p3_add_35454_comb;
  wire [28:0] p3_add_35455_comb;
  wire [31:0] p3_add_35460_comb;
  wire [31:0] p3_add_35461_comb;
  wire [31:0] p3_add_35462_comb;
  wire [31:0] p3_add_35463_comb;
  wire [31:0] p3_add_35464_comb;
  wire [31:0] p3_add_35465_comb;
  wire [31:0] p3_add_35466_comb;
  wire [31:0] p3_add_35467_comb;
  wire [31:0] p3_umul_35468_comb;
  wire [31:0] p3_umul_35469_comb;
  wire [31:0] p3_umul_35470_comb;
  wire [31:0] p3_umul_35471_comb;
  wire [31:0] p3_umul_35472_comb;
  wire [24:0] p3_add_35475_comb;
  wire [20:0] p3_add_35477_comb;
  wire [24:0] p3_add_35481_comb;
  wire [20:0] p3_add_35483_comb;
  wire [24:0] p3_add_35487_comb;
  wire [29:0] p3_add_35488_comb;
  wire [24:0] p3_add_35491_comb;
  wire [28:0] p3_add_35492_comb;
  wire [31:0] p3_sub_35493_comb;
  wire [31:0] p3_sub_35495_comb;
  wire [31:0] p3_sub_35497_comb;
  wire [31:0] p3_sub_35499_comb;
  wire [29:0] p3_add_35511_comb;
  wire [20:0] p3_add_35513_comb;
  wire [28:0] p3_add_35517_comb;
  wire [20:0] p3_add_35519_comb;
  wire [20:0] p3_add_35523_comb;
  wire [20:0] p3_add_35526_comb;
  wire [20:0] p3_add_35531_comb;
  wire [20:0] p3_add_35534_comb;
  wire [31:0] p3_umul_35539_comb;
  wire [31:0] p3_umul_35540_comb;
  wire [31:0] p3_umul_35541_comb;
  wire [31:0] p3_umul_35542_comb;
  wire [29:0] p3_add_35543_comb;
  wire [29:0] p3_add_35546_comb;
  wire [31:0] p3_add_35549_comb;
  wire [31:0] p3_add_35550_comb;
  wire [29:0] p3_add_35551_comb;
  wire [31:0] p3_add_35554_comb;
  wire [31:0] p3_add_35555_comb;
  wire [29:0] p3_add_35556_comb;
  wire [31:0] p3_add_35559_comb;
  wire [31:0] p3_add_35560_comb;
  wire [29:0] p3_add_35561_comb;
  wire [31:0] p3_add_35564_comb;
  wire [31:0] p3_add_35565_comb;
  wire [29:0] p3_add_35573_comb;
  wire [20:0] p3_add_35575_comb;
  wire [28:0] p3_add_35579_comb;
  wire [20:0] p3_add_35581_comb;
  wire [20:0] p3_add_35585_comb;
  wire [20:0] p3_add_35588_comb;
  wire [20:0] p3_add_35593_comb;
  wire [20:0] p3_add_35596_comb;
  wire [31:0] p3_umul_35608_comb;
  wire [31:0] p3_umul_35610_comb;
  wire [31:0] p3_sub_35611_comb;
  wire [31:0] p3_umul_35614_comb;
  wire [31:0] p3_sub_35615_comb;
  wire [31:0] p3_umul_35618_comb;
  wire [31:0] p3_sub_35619_comb;
  wire [31:0] p3_umul_35622_comb;
  wire [31:0] p3_sub_35623_comb;
  wire [31:0] p3_umul_35625_comb;
  wire [31:0] p3_umul_35626_comb;
  wire [31:0] p3_umul_35627_comb;
  wire [31:0] p3_umul_35628_comb;
  wire [31:0] p3_umul_35629_comb;
  wire [31:0] p3_sub_35630_comb;
  wire [31:0] p3_sub_35633_comb;
  wire [31:0] p3_sub_35636_comb;
  wire [31:0] p3_sub_35639_comb;
  wire [24:0] p3_add_35642_comb;
  wire [24:0] p3_add_35643_comb;
  wire [24:0] p3_add_35644_comb;
  wire [24:0] p3_add_35645_comb;
  wire [31:0] p3_sub_35646_comb;
  wire [31:0] p3_sub_35647_comb;
  wire [31:0] p3_umul_35648_comb;
  wire [31:0] p3_sub_35649_comb;
  wire [31:0] p3_umul_35650_comb;
  wire [31:0] p3_sub_35651_comb;
  wire [31:0] p3_umul_35652_comb;
  wire [31:0] p3_sub_35653_comb;
  wire [31:0] p3_umul_35654_comb;
  wire [31:0] p3_sub_35669_comb;
  wire [31:0] p3_sub_35672_comb;
  wire [31:0] p3_sub_35675_comb;
  wire [31:0] p3_sub_35678_comb;
  wire [23:0] p3_bit_slice_35679_comb;
  wire [23:0] p3_bit_slice_35680_comb;
  wire [23:0] p3_bit_slice_35681_comb;
  wire [23:0] p3_bit_slice_35682_comb;
  wire [23:0] p3_bit_slice_35683_comb;
  wire [23:0] p3_bit_slice_35684_comb;
  wire [23:0] p3_bit_slice_35685_comb;
  wire [23:0] p3_bit_slice_35686_comb;
  wire [28:0] p3_bit_slice_35687_comb;
  wire [28:0] p3_bit_slice_35688_comb;
  wire [28:0] p3_bit_slice_35691_comb;
  wire [28:0] p3_bit_slice_35694_comb;
  wire [28:0] p3_bit_slice_35695_comb;
  wire [28:0] p3_bit_slice_35696_comb;
  wire [28:0] p3_bit_slice_35699_comb;
  wire [28:0] p3_bit_slice_35702_comb;
  wire [26:0] p3_add_35703_comb;
  wire [26:0] p3_add_35705_comb;
  wire [26:0] p3_add_35707_comb;
  wire [26:0] p3_add_35709_comb;
  wire [26:0] p3_add_35711_comb;
  wire [18:0] p3_add_35713_comb;
  wire [18:0] p3_add_35718_comb;
  wire [18:0] p3_add_35723_comb;
  wire [18:0] p3_add_35732_comb;
  wire [18:0] p3_add_35737_comb;
  wire [31:0] p3_sign_ext_35744_comb;
  wire [31:0] p3_sign_ext_35745_comb;
  wire [31:0] p3_sign_ext_35746_comb;
  wire [31:0] p3_sign_ext_35747_comb;
  wire [31:0] p3_sign_ext_35748_comb;
  wire [31:0] p3_sign_ext_35749_comb;
  wire [31:0] p3_sign_ext_35750_comb;
  wire [31:0] p3_sign_ext_35751_comb;
  wire [31:0] p3_sign_ext_35752_comb;
  wire [31:0] p3_sign_ext_35753_comb;
  wire [24:0] p3_add_35754_comb;
  wire [31:0] p3_sign_ext_35755_comb;
  wire [24:0] p3_add_35756_comb;
  wire [31:0] p3_sign_ext_35757_comb;
  wire [31:0] p3_sign_ext_35758_comb;
  wire [31:0] p3_sign_ext_35759_comb;
  wire [24:0] p3_add_35760_comb;
  wire [31:0] p3_sign_ext_35761_comb;
  wire [24:0] p3_add_35762_comb;
  wire [31:0] p3_sign_ext_35763_comb;
  wire [28:0] p3_concat_35764_comb;
  wire [28:0] p3_concat_35765_comb;
  wire [28:0] p3_concat_35766_comb;
  wire [28:0] p3_concat_35767_comb;
  wire [28:0] p3_concat_35768_comb;
  wire [31:0] p3_concat_35769_comb;
  wire [31:0] p3_concat_35771_comb;
  wire [31:0] p3_concat_35773_comb;
  wire [31:0] p3_concat_35775_comb;
  wire [31:0] p3_concat_35777_comb;
  wire [31:0] p3_concat_35779_comb;
  wire [31:0] p3_concat_35781_comb;
  wire [31:0] p3_concat_35783_comb;
  wire [23:0] p3_bit_slice_35813_comb;
  wire [23:0] p3_bit_slice_35816_comb;
  wire [23:0] p3_bit_slice_35819_comb;
  wire [23:0] p3_bit_slice_35822_comb;
  wire [23:0] p3_bit_slice_35825_comb;
  wire [23:0] p3_bit_slice_35828_comb;
  wire [23:0] p3_bit_slice_35831_comb;
  wire [23:0] p3_bit_slice_35834_comb;
  wire [31:0] p3_sign_ext_35835_comb;
  wire [31:0] p3_sign_ext_35837_comb;
  wire [31:0] p3_sign_ext_35839_comb;
  wire [31:0] p3_sign_ext_35841_comb;
  wire [31:0] p3_sign_ext_35843_comb;
  wire [31:0] p3_sub_35845_comb;
  wire [31:0] p3_sub_35846_comb;
  wire [31:0] p3_sub_35847_comb;
  wire [31:0] p3_sub_35848_comb;
  wire [31:0] p3_sub_35849_comb;
  wire [31:0] p3_sub_35850_comb;
  wire [31:0] p3_sub_35851_comb;
  wire [31:0] p3_sub_35852_comb;
  wire [18:0] p3_add_35853_comb;
  wire [18:0] p3_add_35855_comb;
  wire [18:0] p3_add_35857_comb;
  wire [18:0] p3_add_35859_comb;
  wire [18:0] p3_add_35861_comb;
  wire [18:0] p3_add_35863_comb;
  wire [18:0] p3_add_35865_comb;
  wire [18:0] p3_add_35867_comb;
  wire [18:0] p3_add_35869_comb;
  wire [18:0] p3_add_35871_comb;
  wire [18:0] p3_add_35873_comb;
  wire [18:0] p3_add_35875_comb;
  wire [18:0] p3_add_35877_comb;
  wire [31:0] p3_add_35879_comb;
  wire [31:0] p3_add_35880_comb;
  wire [31:0] p3_add_35881_comb;
  wire [31:0] p3_add_35882_comb;
  wire [31:0] p3_add_35883_comb;
  wire [31:0] p3_add_35884_comb;
  wire [31:0] p3_add_35885_comb;
  wire [31:0] p3_add_35886_comb;
  wire [18:0] p3_add_35887_comb;
  wire [31:0] p3_sign_ext_35889_comb;
  wire [18:0] p3_add_35890_comb;
  wire [31:0] p3_sign_ext_35892_comb;
  wire [18:0] p3_add_35893_comb;
  wire [31:0] p3_sign_ext_35895_comb;
  wire [18:0] p3_add_35896_comb;
  wire [31:0] p3_sign_ext_35898_comb;
  wire [18:0] p3_add_35899_comb;
  wire [31:0] p3_sign_ext_35901_comb;
  wire [18:0] p3_add_35902_comb;
  wire [31:0] p3_sign_ext_35904_comb;
  wire [18:0] p3_add_35905_comb;
  wire [31:0] p3_sign_ext_35907_comb;
  wire [18:0] p3_add_35908_comb;
  wire [31:0] p3_sign_ext_35910_comb;
  wire [23:0] p3_add_35912_comb;
  wire [23:0] p3_add_35914_comb;
  wire [23:0] p3_add_35916_comb;
  wire [23:0] p3_add_35918_comb;
  wire [23:0] p3_add_35920_comb;
  wire [23:0] p3_add_35984_comb;
  wire [23:0] p3_add_35986_comb;
  wire [23:0] p3_add_35988_comb;
  wire [23:0] p3_add_35990_comb;
  wire [23:0] p3_add_35992_comb;
  wire [23:0] p3_add_35994_comb;
  wire [23:0] p3_add_35996_comb;
  wire [23:0] p3_add_35998_comb;
  wire [23:0] p3_add_36000_comb;
  wire [23:0] p3_add_36002_comb;
  wire [23:0] p3_add_36004_comb;
  wire [23:0] p3_add_36006_comb;
  wire [23:0] p3_add_36008_comb;
  wire [23:0] p3_add_36010_comb;
  wire [23:0] p3_add_36012_comb;
  wire [23:0] p3_add_36013_comb;
  wire [23:0] p3_add_36015_comb;
  wire [23:0] p3_add_36016_comb;
  wire [23:0] p3_add_36018_comb;
  wire [23:0] p3_add_36019_comb;
  wire [23:0] p3_add_36021_comb;
  wire [23:0] p3_add_36022_comb;
  wire [23:0] p3_add_36024_comb;
  wire [23:0] p3_add_36025_comb;
  wire [23:0] p3_add_36027_comb;
  wire [23:0] p3_add_36028_comb;
  wire [23:0] p3_add_36030_comb;
  wire [23:0] p3_add_36031_comb;
  wire [23:0] p3_add_36033_comb;
  wire [23:0] p3_add_36039_comb;
  wire [23:0] p3_add_36041_comb;
  wire [31:0] p3_add_36043_comb;
  wire [23:0] p3_add_36044_comb;
  wire [31:0] p3_add_36046_comb;
  wire [23:0] p3_add_36047_comb;
  wire [31:0] p3_add_36049_comb;
  wire [23:0] p3_add_36050_comb;
  wire [31:0] p3_add_36052_comb;
  wire [23:0] p3_add_36053_comb;
  wire [23:0] p3_add_36055_comb;
  wire [23:0] p3_add_36057_comb;
  wire [23:0] p3_add_36059_comb;
  wire [23:0] p3_add_36061_comb;
  wire [23:0] p3_add_36063_comb;
  wire [23:0] p3_add_36065_comb;
  wire [23:0] p3_add_36067_comb;
  wire [23:0] p3_add_36069_comb;
  wire [23:0] p3_add_36070_comb;
  wire [23:0] p3_add_36072_comb;
  wire [23:0] p3_add_36073_comb;
  wire [23:0] p3_add_36075_comb;
  wire [23:0] p3_add_36076_comb;
  wire [23:0] p3_add_36078_comb;
  wire [23:0] p3_add_36079_comb;
  wire [23:0] p3_add_36081_comb;
  wire [23:0] p3_add_36082_comb;
  wire [23:0] p3_add_36084_comb;
  wire [23:0] p3_add_36085_comb;
  wire [23:0] p3_add_36087_comb;
  wire [23:0] p3_add_36088_comb;
  wire [23:0] p3_add_36090_comb;
  wire [23:0] p3_add_36091_comb;
  wire [31:0] p3_concat_36093_comb;
  wire [31:0] p3_add_36094_comb;
  wire [31:0] p3_concat_36095_comb;
  wire [31:0] p3_add_36096_comb;
  wire [31:0] p3_concat_36097_comb;
  wire [31:0] p3_add_36098_comb;
  wire [31:0] p3_concat_36099_comb;
  wire [31:0] p3_add_36100_comb;
  wire [31:0] p3_concat_36101_comb;
  wire [31:0] p3_sub_36126_comb;
  wire [31:0] p3_sub_36127_comb;
  wire [31:0] p3_sub_36128_comb;
  wire [31:0] p3_sub_36129_comb;
  wire [31:0] p3_sub_36130_comb;
  wire [31:0] p3_add_36132_comb;
  wire [31:0] p3_add_36134_comb;
  wire [31:0] p3_add_36136_comb;
  wire [31:0] p3_add_36138_comb;
  wire [31:0] p3_add_36140_comb;
  wire [31:0] p3_add_36165_comb;
  wire [31:0] p3_add_36166_comb;
  wire [31:0] p3_add_36167_comb;
  wire [31:0] p3_add_36168_comb;
  wire [31:0] p3_add_36169_comb;
  wire [31:0] p3_add_36170_comb;
  wire [31:0] p3_add_36171_comb;
  wire [31:0] p3_add_36172_comb;
  wire [31:0] p3_add_36173_comb;
  wire [31:0] p3_add_36174_comb;
  wire [31:0] p3_add_36175_comb;
  wire [31:0] p3_add_36176_comb;
  wire [31:0] p3_add_36177_comb;
  wire [31:0] p3_sub_36178_comb;
  wire [31:0] p3_sub_36179_comb;
  wire [31:0] p3_sub_36180_comb;
  wire [31:0] p3_sub_36181_comb;
  wire [31:0] p3_sub_36182_comb;
  wire [31:0] p3_sub_36183_comb;
  wire [31:0] p3_sub_36184_comb;
  wire [31:0] p3_sub_36185_comb;
  wire [31:0] p3_add_36186_comb;
  wire [31:0] p3_add_36187_comb;
  wire [31:0] p3_add_36188_comb;
  wire [31:0] p3_add_36189_comb;
  wire [31:0] p3_add_36190_comb;
  wire [31:0] p3_sub_36191_comb;
  wire [31:0] p3_sub_36192_comb;
  wire [31:0] p3_sub_36193_comb;
  wire [31:0] p3_sub_36194_comb;
  wire [31:0] p3_sub_36195_comb;
  wire [31:0] p3_sub_36196_comb;
  wire [31:0] p3_sub_36197_comb;
  wire [31:0] p3_sub_36198_comb;
  wire [31:0] p3_sub_36199_comb;
  wire [31:0] p3_sub_36200_comb;
  wire [31:0] p3_sub_36201_comb;
  wire [31:0] p3_sub_36202_comb;
  wire [31:0] p3_sub_36203_comb;
  wire [31:0] p3_sub_36204_comb;
  wire [31:0] p3_sub_36205_comb;
  wire [31:0] p3_sub_36206_comb;
  wire [31:0] p3_sub_36207_comb;
  wire [31:0] p3_sub_36208_comb;
  wire [31:0] p3_sub_36209_comb;
  wire [31:0] p3_sub_36210_comb;
  wire [31:0] p3_sub_36211_comb;
  wire [31:0] p3_sub_36212_comb;
  wire [31:0] p3_sub_36213_comb;
  wire [31:0] p3_sub_36214_comb;
  wire [31:0] p3_sub_36215_comb;
  wire [31:0] p3_sub_36216_comb;
  wire [17:0] p3_bit_slice_36217_comb;
  wire [17:0] p3_bit_slice_36218_comb;
  wire [17:0] p3_bit_slice_36219_comb;
  wire [17:0] p3_bit_slice_36220_comb;
  wire [17:0] p3_bit_slice_36221_comb;
  wire [17:0] p3_bit_slice_36222_comb;
  wire [17:0] p3_bit_slice_36223_comb;
  wire [17:0] p3_bit_slice_36224_comb;
  wire [17:0] p3_bit_slice_36225_comb;
  wire [17:0] p3_bit_slice_36226_comb;
  wire [17:0] p3_bit_slice_36227_comb;
  wire [17:0] p3_bit_slice_36228_comb;
  wire [17:0] p3_bit_slice_36229_comb;
  wire [17:0] p3_bit_slice_36230_comb;
  wire [17:0] p3_bit_slice_36231_comb;
  wire [17:0] p3_bit_slice_36232_comb;
  wire [17:0] p3_bit_slice_36233_comb;
  wire [17:0] p3_bit_slice_36234_comb;
  wire [17:0] p3_bit_slice_36235_comb;
  wire [17:0] p3_bit_slice_36236_comb;
  wire [17:0] p3_bit_slice_36237_comb;
  wire [17:0] p3_bit_slice_36238_comb;
  wire [17:0] p3_bit_slice_36239_comb;
  wire [17:0] p3_bit_slice_36240_comb;
  wire [17:0] p3_bit_slice_36241_comb;
  wire [17:0] p3_bit_slice_36242_comb;
  wire [17:0] p3_bit_slice_36243_comb;
  wire [17:0] p3_bit_slice_36244_comb;
  wire [17:0] p3_bit_slice_36245_comb;
  wire [17:0] p3_bit_slice_36246_comb;
  wire [17:0] p3_bit_slice_36247_comb;
  wire [17:0] p3_bit_slice_36248_comb;
  wire [17:0] p3_bit_slice_36249_comb;
  wire [17:0] p3_bit_slice_36250_comb;
  wire [17:0] p3_bit_slice_36251_comb;
  wire [17:0] p3_bit_slice_36252_comb;
  wire [17:0] p3_bit_slice_36253_comb;
  wire [17:0] p3_bit_slice_36254_comb;
  wire [17:0] p3_bit_slice_36255_comb;
  wire [17:0] p3_bit_slice_36256_comb;
  wire [17:0] p3_bit_slice_36257_comb;
  wire [17:0] p3_bit_slice_36258_comb;
  wire [17:0] p3_bit_slice_36259_comb;
  wire [17:0] p3_bit_slice_36260_comb;
  wire [17:0] p3_bit_slice_36261_comb;
  wire [17:0] p3_bit_slice_36262_comb;
  wire [17:0] p3_bit_slice_36263_comb;
  wire [17:0] p3_bit_slice_36264_comb;
  wire [17:0] p3_bit_slice_36265_comb;
  wire [17:0] p3_bit_slice_36266_comb;
  wire [17:0] p3_bit_slice_36267_comb;
  wire [17:0] p3_bit_slice_36268_comb;
  wire [31:0] p3_array_36333_comb[64];
  assign p3_bit_slice_35376_comb = p2_add_34680[24:1];
  assign p3_bit_slice_35377_comb = p2_add_34683[24:1];
  assign p3_sign_ext_35378_comb = {{8{p3_bit_slice_35376_comb[23]}}, p3_bit_slice_35376_comb};
  assign p3_bit_slice_35379_comb = p2_add_34747[24:1];
  assign p3_sign_ext_35380_comb = {{8{p3_bit_slice_35377_comb[23]}}, p3_bit_slice_35377_comb};
  assign p3_bit_slice_35381_comb = p2_add_34749[24:1];
  assign p3_sign_ext_35382_comb = {{8{p2_bit_slice_33771[23]}}, p2_bit_slice_33771};
  assign p3_sign_ext_35383_comb = {{8{p2_bit_slice_33772[23]}}, p2_bit_slice_33772};
  assign p3_sign_ext_35384_comb = {{8{p2_bit_slice_34786[23]}}, p2_bit_slice_34786};
  assign p3_sign_ext_35385_comb = {{8{p2_bit_slice_34787[23]}}, p2_bit_slice_34787};
  assign p3_sign_ext_35386_comb = {{8{p2_bit_slice_34788[23]}}, p2_bit_slice_34788};
  assign p3_sign_ext_35387_comb = {{8{p2_bit_slice_34789[23]}}, p2_bit_slice_34789};
  assign p3_sign_ext_35388_comb = {{8{p2_bit_slice_34790[23]}}, p2_bit_slice_34790};
  assign p3_sign_ext_35389_comb = {{8{p2_bit_slice_34791[23]}}, p2_bit_slice_34791};
  assign p3_sign_ext_35390_comb = {{8{p2_bit_slice_34792[23]}}, p2_bit_slice_34792};
  assign p3_sign_ext_35391_comb = {{8{p2_bit_slice_34793[23]}}, p2_bit_slice_34793};
  assign p3_sign_ext_35395_comb = {{8{p3_bit_slice_35379_comb[23]}}, p3_bit_slice_35379_comb};
  assign p3_sign_ext_35399_comb = {{8{p3_bit_slice_35381_comb[23]}}, p3_bit_slice_35381_comb};
  assign p3_sign_ext_35408_comb = {{3{p2_bit_slice_34803[28]}}, p2_bit_slice_34803};
  assign p3_sign_ext_35409_comb = {{3{p2_bit_slice_34804[28]}}, p2_bit_slice_34804};
  assign p3_sign_ext_35410_comb = {{3{p2_bit_slice_34805[28]}}, p2_bit_slice_34805};
  assign p3_sign_ext_35411_comb = {{3{p2_bit_slice_34806[28]}}, p2_bit_slice_34806};
  assign p3_sign_ext_35412_comb = {{3{p2_bit_slice_34807[28]}}, p2_bit_slice_34807};
  assign p3_sign_ext_35413_comb = {{3{p2_bit_slice_34808[28]}}, p2_bit_slice_34808};
  assign p3_sign_ext_35414_comb = {{3{p2_bit_slice_34809[28]}}, p2_bit_slice_34809};
  assign p3_sign_ext_35415_comb = {{3{p2_bit_slice_34810[28]}}, p2_bit_slice_34810};
  assign p3_sign_ext_35416_comb = {{3{p2_bit_slice_34819[28]}}, p2_bit_slice_34819};
  assign p3_sign_ext_35417_comb = {{3{p2_bit_slice_34820[28]}}, p2_bit_slice_34820};
  assign p3_sign_ext_35418_comb = {{3{p2_bit_slice_34821[28]}}, p2_bit_slice_34821};
  assign p3_sign_ext_35419_comb = {{3{p2_bit_slice_34822[28]}}, p2_bit_slice_34822};
  assign p3_sign_ext_35420_comb = {{3{p2_bit_slice_34823[28]}}, p2_bit_slice_34823};
  assign p3_sign_ext_35421_comb = {{3{p2_bit_slice_34824[28]}}, p2_bit_slice_34824};
  assign p3_sign_ext_35422_comb = {{3{p2_bit_slice_34825[28]}}, p2_bit_slice_34825};
  assign p3_sign_ext_35423_comb = {{3{p2_bit_slice_34826[28]}}, p2_bit_slice_34826};
  assign p3_add_35424_comb = p3_sign_ext_35382_comb + p3_sign_ext_35383_comb;
  assign p3_add_35426_comb = p3_sign_ext_35384_comb + p3_sign_ext_35385_comb;
  assign p3_add_35428_comb = p3_sign_ext_35386_comb + p3_sign_ext_35387_comb;
  assign p3_add_35430_comb = p3_sign_ext_35388_comb + p3_sign_ext_35389_comb;
  assign p3_add_35432_comb = p3_sign_ext_35390_comb + p3_sign_ext_35391_comb;
  assign p3_add_35434_comb = p3_sign_ext_35378_comb[31:7] + 25'h000_0001;
  assign p3_add_35436_comb = p2_umul_34687[31:11] + p2_bit_slice_33780;
  assign p3_add_35441_comb = p3_sign_ext_35380_comb[31:7] + 25'h000_0001;
  assign p3_add_35443_comb = p2_umul_34794[31:11] + p2_bit_slice_33780;
  assign p3_add_35448_comb = p2_umul_34794[31:7] + 25'h000_0001;
  assign p3_add_35449_comb = p3_sign_ext_35380_comb[31:2] + p2_umul_34687[31:2];
  assign p3_add_35454_comb = p2_umul_34687[31:7] + 25'h000_0001;
  assign p3_add_35455_comb = p3_sign_ext_35378_comb[31:3] + p2_umul_34794[31:3];
  assign p3_add_35460_comb = p3_sign_ext_35408_comb + p3_sign_ext_35409_comb;
  assign p3_add_35461_comb = p3_sign_ext_35410_comb + p3_sign_ext_35411_comb;
  assign p3_add_35462_comb = p3_sign_ext_35412_comb + p3_sign_ext_35413_comb;
  assign p3_add_35463_comb = p3_sign_ext_35414_comb + p3_sign_ext_35415_comb;
  assign p3_add_35464_comb = p3_sign_ext_35416_comb + p3_sign_ext_35417_comb;
  assign p3_add_35465_comb = p3_sign_ext_35418_comb + p3_sign_ext_35419_comb;
  assign p3_add_35466_comb = p3_sign_ext_35420_comb + p3_sign_ext_35421_comb;
  assign p3_add_35467_comb = p3_sign_ext_35422_comb + p3_sign_ext_35423_comb;
  assign p3_umul_35468_comb = umul32b_32b_x_11b(p3_add_35424_comb, 11'h454);
  assign p3_umul_35469_comb = umul32b_32b_x_11b(p3_add_35426_comb, 11'h454);
  assign p3_umul_35470_comb = umul32b_32b_x_11b(p3_add_35428_comb, 11'h454);
  assign p3_umul_35471_comb = umul32b_32b_x_11b(p3_add_35430_comb, 11'h454);
  assign p3_umul_35472_comb = umul32b_32b_x_11b(p3_add_35432_comb, 11'h454);
  assign p3_add_35475_comb = p3_sign_ext_35395_comb[31:7] + 25'h000_0001;
  assign p3_add_35477_comb = p2_umul_34753[31:11] + p2_bit_slice_33784;
  assign p3_add_35481_comb = p3_sign_ext_35399_comb[31:7] + 25'h000_0001;
  assign p3_add_35483_comb = p2_umul_34837[31:11] + p2_bit_slice_33784;
  assign p3_add_35487_comb = p2_umul_34837[31:7] + 25'h000_0001;
  assign p3_add_35488_comb = p3_sign_ext_35399_comb[31:2] + p2_umul_34753[31:2];
  assign p3_add_35491_comb = p2_umul_34753[31:7] + 25'h000_0001;
  assign p3_add_35492_comb = p3_sign_ext_35395_comb[31:3] + p2_umul_34837[31:3];
  assign p3_sub_35493_comb = p3_add_35460_comb - p3_add_35461_comb;
  assign p3_sub_35495_comb = p3_add_35462_comb - p3_add_35463_comb;
  assign p3_sub_35497_comb = p3_add_35464_comb - p3_add_35465_comb;
  assign p3_sub_35499_comb = p3_add_35466_comb - p3_add_35467_comb;
  assign p3_add_35511_comb = {p3_add_35434_comb, p2_add_34680[7:3]} + {p3_add_35436_comb, p2_umul_34687[10:2]};
  assign p3_add_35513_comb = p2_umul_34794[31:11] + p2_bit_slice_33779;
  assign p3_add_35517_comb = {p3_add_35441_comb, p2_add_34683[7:4]} + {p3_add_35443_comb, p2_umul_34794[10:3]};
  assign p3_add_35519_comb = p2_umul_34687[31:11] + p2_bit_slice_33779;
  assign p3_add_35523_comb = p3_add_35448_comb[24:4] + p2_bit_slice_33780;
  assign p3_add_35526_comb = p3_add_35449_comb[29:9] + p2_bit_slice_33779;
  assign p3_add_35531_comb = p3_add_35454_comb[24:4] + p2_bit_slice_33780;
  assign p3_add_35534_comb = p3_add_35455_comb[28:8] + p2_bit_slice_33779;
  assign p3_umul_35539_comb = umul32b_32b_x_8b(p3_sub_35493_comb, 8'hb5);
  assign p3_umul_35540_comb = umul32b_32b_x_8b(p3_sub_35495_comb, 8'hb5);
  assign p3_umul_35541_comb = umul32b_32b_x_8b(p3_sub_35497_comb, 8'hb5);
  assign p3_umul_35542_comb = umul32b_32b_x_8b(p3_sub_35499_comb, 8'hb5);
  assign p3_add_35543_comb = p3_umul_35468_comb[31:2] + 30'h0000_0001;
  assign p3_add_35546_comb = p3_umul_35469_comb[31:2] + 30'h0000_0001;
  assign p3_add_35549_comb = p3_sign_ext_35408_comb + p3_sign_ext_35411_comb;
  assign p3_add_35550_comb = p3_sign_ext_35410_comb + p3_sign_ext_35409_comb;
  assign p3_add_35551_comb = p3_umul_35470_comb[31:2] + 30'h0000_0001;
  assign p3_add_35554_comb = p3_sign_ext_35412_comb + p3_sign_ext_35415_comb;
  assign p3_add_35555_comb = p3_sign_ext_35414_comb + p3_sign_ext_35413_comb;
  assign p3_add_35556_comb = p3_umul_35471_comb[31:2] + 30'h0000_0001;
  assign p3_add_35559_comb = p3_sign_ext_35416_comb + p3_sign_ext_35419_comb;
  assign p3_add_35560_comb = p3_sign_ext_35418_comb + p3_sign_ext_35417_comb;
  assign p3_add_35561_comb = p3_umul_35472_comb[31:2] + 30'h0000_0001;
  assign p3_add_35564_comb = p3_sign_ext_35420_comb + p3_sign_ext_35423_comb;
  assign p3_add_35565_comb = p3_sign_ext_35422_comb + p3_sign_ext_35421_comb;
  assign p3_add_35573_comb = {p3_add_35475_comb, p2_add_34747[7:3]} + {p3_add_35477_comb, p2_umul_34753[10:2]};
  assign p3_add_35575_comb = p2_umul_34837[31:11] + p2_bit_slice_33783;
  assign p3_add_35579_comb = {p3_add_35481_comb, p2_add_34749[7:4]} + {p3_add_35483_comb, p2_umul_34837[10:3]};
  assign p3_add_35581_comb = p2_umul_34753[31:11] + p2_bit_slice_33783;
  assign p3_add_35585_comb = p3_add_35487_comb[24:4] + p2_bit_slice_33784;
  assign p3_add_35588_comb = p3_add_35488_comb[29:9] + p2_bit_slice_33783;
  assign p3_add_35593_comb = p3_add_35491_comb[24:4] + p2_bit_slice_33784;
  assign p3_add_35596_comb = p3_add_35492_comb[28:8] + p2_bit_slice_33783;
  assign p3_umul_35608_comb = umul32b_32b_x_12b(p3_sign_ext_35383_comb, 12'hec8);
  assign p3_umul_35610_comb = umul32b_32b_x_12b(p3_sign_ext_35385_comb, 12'hec8);
  assign p3_sub_35611_comb = p3_add_35549_comb - p3_add_35550_comb;
  assign p3_umul_35614_comb = umul32b_32b_x_12b(p3_sign_ext_35387_comb, 12'hec8);
  assign p3_sub_35615_comb = p3_add_35554_comb - p3_add_35555_comb;
  assign p3_umul_35618_comb = umul32b_32b_x_12b(p3_sign_ext_35389_comb, 12'hec8);
  assign p3_sub_35619_comb = p3_add_35559_comb - p3_add_35560_comb;
  assign p3_umul_35622_comb = umul32b_32b_x_12b(p3_sign_ext_35391_comb, 12'hec8);
  assign p3_sub_35623_comb = p3_add_35564_comb - p3_add_35565_comb;
  assign p3_umul_35625_comb = umul32b_32b_x_11b(p3_sign_ext_35382_comb, 11'h620);
  assign p3_umul_35626_comb = umul32b_32b_x_11b(p3_sign_ext_35384_comb, 11'h620);
  assign p3_umul_35627_comb = umul32b_32b_x_11b(p3_sign_ext_35386_comb, 11'h620);
  assign p3_umul_35628_comb = umul32b_32b_x_11b(p3_sign_ext_35388_comb, 11'h620);
  assign p3_umul_35629_comb = umul32b_32b_x_11b(p3_sign_ext_35390_comb, 11'h620);
  assign p3_sub_35630_comb = {p3_add_35511_comb, p2_add_34680[2:1]} - {p3_add_35513_comb, p2_umul_34794[10:0]};
  assign p3_sub_35633_comb = {p3_add_35517_comb, p2_add_34683[3:1]} - {p3_add_35519_comb, p2_umul_34687[10:0]};
  assign p3_sub_35636_comb = {p3_add_35523_comb, p3_add_35448_comb[3:0], p2_umul_34794[6:0]} - {p3_add_35526_comb, p3_add_35449_comb[8:0], p2_add_34683[2:1]};
  assign p3_sub_35639_comb = {p3_add_35531_comb, p3_add_35454_comb[3:0], p2_umul_34687[6:0]} - {p3_add_35534_comb, p3_add_35455_comb[7:0], p2_add_34680[3:1]};
  assign p3_add_35642_comb = p3_umul_35539_comb[31:7] + 25'h000_0001;
  assign p3_add_35643_comb = p3_umul_35540_comb[31:7] + 25'h000_0001;
  assign p3_add_35644_comb = p3_umul_35541_comb[31:7] + 25'h000_0001;
  assign p3_add_35645_comb = p3_umul_35542_comb[31:7] + 25'h000_0001;
  assign p3_sub_35646_comb = {p3_add_35543_comb, 2'h0} - p3_umul_35608_comb;
  assign p3_sub_35647_comb = {p3_add_35546_comb, 2'h0} - p3_umul_35610_comb;
  assign p3_umul_35648_comb = umul32b_32b_x_8b(p3_sub_35611_comb, 8'hb5);
  assign p3_sub_35649_comb = {p3_add_35551_comb, 2'h0} - p3_umul_35614_comb;
  assign p3_umul_35650_comb = umul32b_32b_x_8b(p3_sub_35615_comb, 8'hb5);
  assign p3_sub_35651_comb = {p3_add_35556_comb, 2'h0} - p3_umul_35618_comb;
  assign p3_umul_35652_comb = umul32b_32b_x_8b(p3_sub_35619_comb, 8'hb5);
  assign p3_sub_35653_comb = {p3_add_35561_comb, 2'h0} - p3_umul_35622_comb;
  assign p3_umul_35654_comb = umul32b_32b_x_8b(p3_sub_35623_comb, 8'hb5);
  assign p3_sub_35669_comb = {p3_add_35573_comb, p2_add_34747[2:1]} - {p3_add_35575_comb, p2_umul_34837[10:0]};
  assign p3_sub_35672_comb = {p3_add_35579_comb, p2_add_34749[3:1]} - {p3_add_35581_comb, p2_umul_34753[10:0]};
  assign p3_sub_35675_comb = {p3_add_35585_comb, p3_add_35487_comb[3:0], p2_umul_34837[6:0]} - {p3_add_35588_comb, p3_add_35488_comb[8:0], p2_add_34749[2:1]};
  assign p3_sub_35678_comb = {p3_add_35593_comb, p3_add_35491_comb[3:0], p2_umul_34753[6:0]} - {p3_add_35596_comb, p3_add_35492_comb[7:0], p2_add_34747[3:1]};
  assign p3_bit_slice_35679_comb = p2_add_35073[24:1];
  assign p3_bit_slice_35680_comb = p3_add_35642_comb[24:1];
  assign p3_bit_slice_35681_comb = p3_add_35643_comb[24:1];
  assign p3_bit_slice_35682_comb = p2_add_35074[24:1];
  assign p3_bit_slice_35683_comb = p2_add_35075[24:1];
  assign p3_bit_slice_35684_comb = p3_add_35644_comb[24:1];
  assign p3_bit_slice_35685_comb = p3_add_35645_comb[24:1];
  assign p3_bit_slice_35686_comb = p2_add_35076[24:1];
  assign p3_bit_slice_35687_comb = p3_sub_35646_comb[31:3];
  assign p3_bit_slice_35688_comb = p3_sub_35647_comb[31:3];
  assign p3_bit_slice_35691_comb = p3_sub_35649_comb[31:3];
  assign p3_bit_slice_35694_comb = p2_sub_35078[31:3];
  assign p3_bit_slice_35695_comb = p2_sub_35080[31:3];
  assign p3_bit_slice_35696_comb = p3_sub_35651_comb[31:3];
  assign p3_bit_slice_35699_comb = p3_sub_35653_comb[31:3];
  assign p3_bit_slice_35702_comb = p2_sub_35082[31:3];
  assign p3_add_35703_comb = p3_umul_35625_comb[31:5] + p3_add_35543_comb[29:3];
  assign p3_add_35705_comb = p3_umul_35626_comb[31:5] + p3_add_35546_comb[29:3];
  assign p3_add_35707_comb = p3_umul_35627_comb[31:5] + p3_add_35551_comb[29:3];
  assign p3_add_35709_comb = p3_umul_35628_comb[31:5] + p3_add_35556_comb[29:3];
  assign p3_add_35711_comb = p3_umul_35629_comb[31:5] + p3_add_35561_comb[29:3];
  assign p3_add_35713_comb = p2_add_35061[29:11] + 19'h0_0001;
  assign p3_add_35718_comb = p3_sub_35630_comb[31:13] + 19'h0_0001;
  assign p3_add_35723_comb = p3_sub_35633_comb[31:13] + 19'h0_0001;
  assign p3_add_35732_comb = p3_sub_35636_comb[31:13] + 19'h0_0001;
  assign p3_add_35737_comb = p3_sub_35639_comb[31:13] + 19'h0_0001;
  assign p3_sign_ext_35744_comb = {{8{p3_bit_slice_35679_comb[23]}}, p3_bit_slice_35679_comb};
  assign p3_sign_ext_35745_comb = {{8{p3_bit_slice_35680_comb[23]}}, p3_bit_slice_35680_comb};
  assign p3_sign_ext_35746_comb = {{8{p3_bit_slice_35681_comb[23]}}, p3_bit_slice_35681_comb};
  assign p3_sign_ext_35747_comb = {{8{p3_bit_slice_35682_comb[23]}}, p3_bit_slice_35682_comb};
  assign p3_sign_ext_35748_comb = {{8{p3_bit_slice_35683_comb[23]}}, p3_bit_slice_35683_comb};
  assign p3_sign_ext_35749_comb = {{8{p3_bit_slice_35684_comb[23]}}, p3_bit_slice_35684_comb};
  assign p3_sign_ext_35750_comb = {{8{p3_bit_slice_35685_comb[23]}}, p3_bit_slice_35685_comb};
  assign p3_sign_ext_35751_comb = {{8{p3_bit_slice_35686_comb[23]}}, p3_bit_slice_35686_comb};
  assign p3_sign_ext_35752_comb = {{3{p3_bit_slice_35687_comb[28]}}, p3_bit_slice_35687_comb};
  assign p3_sign_ext_35753_comb = {{3{p3_bit_slice_35688_comb[28]}}, p3_bit_slice_35688_comb};
  assign p3_add_35754_comb = p3_umul_35648_comb[31:7] + 25'h000_0001;
  assign p3_sign_ext_35755_comb = {{3{p3_bit_slice_35691_comb[28]}}, p3_bit_slice_35691_comb};
  assign p3_add_35756_comb = p3_umul_35650_comb[31:7] + 25'h000_0001;
  assign p3_sign_ext_35757_comb = {{3{p3_bit_slice_35694_comb[28]}}, p3_bit_slice_35694_comb};
  assign p3_sign_ext_35758_comb = {{3{p3_bit_slice_35695_comb[28]}}, p3_bit_slice_35695_comb};
  assign p3_sign_ext_35759_comb = {{3{p3_bit_slice_35696_comb[28]}}, p3_bit_slice_35696_comb};
  assign p3_add_35760_comb = p3_umul_35652_comb[31:7] + 25'h000_0001;
  assign p3_sign_ext_35761_comb = {{3{p3_bit_slice_35699_comb[28]}}, p3_bit_slice_35699_comb};
  assign p3_add_35762_comb = p3_umul_35654_comb[31:7] + 25'h000_0001;
  assign p3_sign_ext_35763_comb = {{3{p3_bit_slice_35702_comb[28]}}, p3_bit_slice_35702_comb};
  assign p3_concat_35764_comb = {p3_add_35703_comb, p3_add_35543_comb[2:1]};
  assign p3_concat_35765_comb = {p3_add_35705_comb, p3_add_35546_comb[2:1]};
  assign p3_concat_35766_comb = {p3_add_35707_comb, p3_add_35551_comb[2:1]};
  assign p3_concat_35767_comb = {p3_add_35709_comb, p3_add_35556_comb[2:1]};
  assign p3_concat_35768_comb = {p3_add_35711_comb, p3_add_35561_comb[2:1]};
  assign p3_concat_35769_comb = {p3_add_35713_comb, p2_add_35061[10:6], 8'h00};
  assign p3_concat_35771_comb = {p3_add_35718_comb, p3_sub_35630_comb[12:8], 8'h00};
  assign p3_concat_35773_comb = {p3_add_35723_comb, p3_sub_35633_comb[12:8], 8'h00};
  assign p3_concat_35775_comb = {p2_add_35114, p2_bit_slice_35115, 8'h00};
  assign p3_concat_35777_comb = {p2_add_35117, p2_bit_slice_35118, 8'h00};
  assign p3_concat_35779_comb = {p3_add_35732_comb, p3_sub_35636_comb[12:8], 8'h00};
  assign p3_concat_35781_comb = {p3_add_35737_comb, p3_sub_35639_comb[12:8], 8'h00};
  assign p3_concat_35783_comb = {p2_add_35120, p2_bit_slice_35121, 8'h00};
  assign p3_bit_slice_35813_comb = p2_add_35123[24:1];
  assign p3_bit_slice_35816_comb = p3_add_35754_comb[24:1];
  assign p3_bit_slice_35819_comb = p3_add_35756_comb[24:1];
  assign p3_bit_slice_35822_comb = p2_add_35124[24:1];
  assign p3_bit_slice_35825_comb = p2_add_35125[24:1];
  assign p3_bit_slice_35828_comb = p3_add_35760_comb[24:1];
  assign p3_bit_slice_35831_comb = p3_add_35762_comb[24:1];
  assign p3_bit_slice_35834_comb = p2_add_35126[24:1];
  assign p3_sign_ext_35835_comb = {{3{p3_concat_35764_comb[28]}}, p3_concat_35764_comb};
  assign p3_sign_ext_35837_comb = {{3{p3_concat_35765_comb[28]}}, p3_concat_35765_comb};
  assign p3_sign_ext_35839_comb = {{3{p3_concat_35766_comb[28]}}, p3_concat_35766_comb};
  assign p3_sign_ext_35841_comb = {{3{p3_concat_35767_comb[28]}}, p3_concat_35767_comb};
  assign p3_sign_ext_35843_comb = {{3{p3_concat_35768_comb[28]}}, p3_concat_35768_comb};
  assign p3_sub_35845_comb = p3_concat_35769_comb - {p2_add_35090[29:6], 8'h00};
  assign p3_sub_35846_comb = p3_concat_35771_comb - {p3_sub_35669_comb[31:8], 8'h00};
  assign p3_sub_35847_comb = p3_concat_35773_comb - {p3_sub_35672_comb[31:8], 8'h00};
  assign p3_sub_35848_comb = p3_concat_35775_comb - {p2_bit_slice_35116, 8'h00};
  assign p3_sub_35849_comb = p3_concat_35777_comb - {p2_bit_slice_35119, 8'h00};
  assign p3_sub_35850_comb = p3_concat_35779_comb - {p3_sub_35675_comb[31:8], 8'h00};
  assign p3_sub_35851_comb = p3_concat_35781_comb - {p3_sub_35678_comb[31:8], 8'h00};
  assign p3_sub_35852_comb = p3_concat_35783_comb - {p2_bit_slice_35122, 8'h00};
  assign p3_add_35853_comb = p3_sign_ext_35744_comb[31:13] + 19'h0_0001;
  assign p3_add_35855_comb = p3_sign_ext_35745_comb[31:13] + 19'h0_0001;
  assign p3_add_35857_comb = p3_sign_ext_35746_comb[31:13] + 19'h0_0001;
  assign p3_add_35859_comb = p3_sign_ext_35747_comb[31:13] + 19'h0_0001;
  assign p3_add_35861_comb = p3_sign_ext_35748_comb[31:13] + 19'h0_0001;
  assign p3_add_35863_comb = p3_sign_ext_35749_comb[31:13] + 19'h0_0001;
  assign p3_add_35865_comb = p3_sign_ext_35750_comb[31:13] + 19'h0_0001;
  assign p3_add_35867_comb = p3_sign_ext_35751_comb[31:13] + 19'h0_0001;
  assign p3_add_35869_comb = p2_add_35090[29:11] + 19'h0_0001;
  assign p3_add_35871_comb = p3_sub_35669_comb[31:13] + 19'h0_0001;
  assign p3_add_35873_comb = p3_sub_35672_comb[31:13] + 19'h0_0001;
  assign p3_add_35875_comb = p3_sub_35675_comb[31:13] + 19'h0_0001;
  assign p3_add_35877_comb = p3_sub_35678_comb[31:13] + 19'h0_0001;
  assign p3_add_35879_comb = p3_sign_ext_35744_comb + p3_sign_ext_35752_comb;
  assign p3_add_35880_comb = p3_sign_ext_35745_comb + p3_sign_ext_35753_comb;
  assign p3_add_35881_comb = p3_sign_ext_35746_comb + p3_sign_ext_35755_comb;
  assign p3_add_35882_comb = p3_sign_ext_35747_comb + p3_sign_ext_35757_comb;
  assign p3_add_35883_comb = p3_sign_ext_35748_comb + p3_sign_ext_35758_comb;
  assign p3_add_35884_comb = p3_sign_ext_35749_comb + p3_sign_ext_35759_comb;
  assign p3_add_35885_comb = p3_sign_ext_35750_comb + p3_sign_ext_35761_comb;
  assign p3_add_35886_comb = p3_sign_ext_35751_comb + p3_sign_ext_35763_comb;
  assign p3_add_35887_comb = p3_sign_ext_35752_comb[31:13] + 19'h0_0001;
  assign p3_sign_ext_35889_comb = {{8{p3_bit_slice_35813_comb[23]}}, p3_bit_slice_35813_comb};
  assign p3_add_35890_comb = p3_sign_ext_35753_comb[31:13] + 19'h0_0001;
  assign p3_sign_ext_35892_comb = {{8{p3_bit_slice_35816_comb[23]}}, p3_bit_slice_35816_comb};
  assign p3_add_35893_comb = p3_sign_ext_35755_comb[31:13] + 19'h0_0001;
  assign p3_sign_ext_35895_comb = {{8{p3_bit_slice_35819_comb[23]}}, p3_bit_slice_35819_comb};
  assign p3_add_35896_comb = p3_sign_ext_35757_comb[31:13] + 19'h0_0001;
  assign p3_sign_ext_35898_comb = {{8{p3_bit_slice_35822_comb[23]}}, p3_bit_slice_35822_comb};
  assign p3_add_35899_comb = p3_sign_ext_35758_comb[31:13] + 19'h0_0001;
  assign p3_sign_ext_35901_comb = {{8{p3_bit_slice_35825_comb[23]}}, p3_bit_slice_35825_comb};
  assign p3_add_35902_comb = p3_sign_ext_35759_comb[31:13] + 19'h0_0001;
  assign p3_sign_ext_35904_comb = {{8{p3_bit_slice_35828_comb[23]}}, p3_bit_slice_35828_comb};
  assign p3_add_35905_comb = p3_sign_ext_35761_comb[31:13] + 19'h0_0001;
  assign p3_sign_ext_35907_comb = {{8{p3_bit_slice_35831_comb[23]}}, p3_bit_slice_35831_comb};
  assign p3_add_35908_comb = p3_sign_ext_35763_comb[31:13] + 19'h0_0001;
  assign p3_sign_ext_35910_comb = {{8{p3_bit_slice_35834_comb[23]}}, p3_bit_slice_35834_comb};
  assign p3_add_35912_comb = p2_add_35090[29:6] + {p3_add_35713_comb, p2_add_35061[10:6]};
  assign p3_add_35914_comb = p3_sub_35669_comb[31:8] + {p3_add_35718_comb, p3_sub_35630_comb[12:8]};
  assign p3_add_35916_comb = p3_sub_35672_comb[31:8] + {p3_add_35723_comb, p3_sub_35633_comb[12:8]};
  assign p3_add_35918_comb = p3_sub_35675_comb[31:8] + {p3_add_35732_comb, p3_sub_35636_comb[12:8]};
  assign p3_add_35920_comb = p3_sub_35678_comb[31:8] + {p3_add_35737_comb, p3_sub_35639_comb[12:8]};
  assign p3_add_35984_comb = p3_sign_ext_35835_comb[31:8] + p3_add_35912_comb;
  assign p3_add_35986_comb = p3_sign_ext_35837_comb[31:8] + p3_add_35914_comb;
  assign p3_add_35988_comb = p3_sign_ext_35839_comb[31:8] + p3_add_35916_comb;
  assign p3_add_35990_comb = p3_sign_ext_35841_comb[31:8] + p3_add_35918_comb;
  assign p3_add_35992_comb = p3_sign_ext_35843_comb[31:8] + p3_add_35920_comb;
  assign p3_add_35994_comb = p3_sign_ext_35752_comb[31:8] + p3_sub_35845_comb[31:8];
  assign p3_add_35996_comb = p3_sign_ext_35753_comb[31:8] + p3_sub_35846_comb[31:8];
  assign p3_add_35998_comb = p3_sign_ext_35755_comb[31:8] + p3_sub_35847_comb[31:8];
  assign p3_add_36000_comb = p3_sign_ext_35757_comb[31:8] + p3_sub_35848_comb[31:8];
  assign p3_add_36002_comb = p3_sign_ext_35758_comb[31:8] + p3_sub_35849_comb[31:8];
  assign p3_add_36004_comb = p3_sign_ext_35759_comb[31:8] + p3_sub_35850_comb[31:8];
  assign p3_add_36006_comb = p3_sign_ext_35761_comb[31:8] + p3_sub_35851_comb[31:8];
  assign p3_add_36008_comb = p3_sign_ext_35763_comb[31:8] + p3_sub_35852_comb[31:8];
  assign p3_add_36010_comb = {p3_add_35853_comb, p2_add_35073[13:9]} + p2_add_35061[29:6];
  assign p3_add_36012_comb = p3_sign_ext_35752_comb[31:8] + p2_add_35090[29:6];
  assign p3_add_36013_comb = {p3_add_35855_comb, p3_add_35642_comb[13:9]} + p3_sub_35630_comb[31:8];
  assign p3_add_36015_comb = p3_sign_ext_35753_comb[31:8] + p3_sub_35669_comb[31:8];
  assign p3_add_36016_comb = {p3_add_35857_comb, p3_add_35643_comb[13:9]} + p3_sub_35633_comb[31:8];
  assign p3_add_36018_comb = p3_sign_ext_35755_comb[31:8] + p3_sub_35672_comb[31:8];
  assign p3_add_36019_comb = {p3_add_35859_comb, p2_add_35074[13:9]} + p2_bit_slice_35154;
  assign p3_add_36021_comb = p3_sign_ext_35757_comb[31:8] + p2_bit_slice_35116;
  assign p3_add_36022_comb = {p3_add_35861_comb, p2_add_35075[13:9]} + p2_bit_slice_35155;
  assign p3_add_36024_comb = p3_sign_ext_35758_comb[31:8] + p2_bit_slice_35119;
  assign p3_add_36025_comb = {p3_add_35863_comb, p3_add_35644_comb[13:9]} + p3_sub_35636_comb[31:8];
  assign p3_add_36027_comb = p3_sign_ext_35759_comb[31:8] + p3_sub_35675_comb[31:8];
  assign p3_add_36028_comb = {p3_add_35865_comb, p3_add_35645_comb[13:9]} + p3_sub_35639_comb[31:8];
  assign p3_add_36030_comb = p3_sign_ext_35761_comb[31:8] + p3_sub_35678_comb[31:8];
  assign p3_add_36031_comb = {p3_add_35867_comb, p2_add_35076[13:9]} + p2_bit_slice_35156;
  assign p3_add_36033_comb = p3_sign_ext_35763_comb[31:8] + p2_bit_slice_35122;
  assign p3_add_36039_comb = {p3_add_35869_comb, p2_add_35090[10:6]} + p2_add_35061[29:6];
  assign p3_add_36041_comb = {p3_add_35871_comb, p3_sub_35669_comb[12:8]} + p3_sub_35630_comb[31:8];
  assign p3_add_36043_comb = p3_sign_ext_35409_comb + p3_sign_ext_35411_comb;
  assign p3_add_36044_comb = {p3_add_35873_comb, p3_sub_35672_comb[12:8]} + p3_sub_35633_comb[31:8];
  assign p3_add_36046_comb = p3_sign_ext_35413_comb + p3_sign_ext_35415_comb;
  assign p3_add_36047_comb = {p3_add_35875_comb, p3_sub_35675_comb[12:8]} + p3_sub_35636_comb[31:8];
  assign p3_add_36049_comb = p3_sign_ext_35417_comb + p3_sign_ext_35419_comb;
  assign p3_add_36050_comb = {p3_add_35877_comb, p3_sub_35678_comb[12:8]} + p3_sub_35639_comb[31:8];
  assign p3_add_36052_comb = p3_sign_ext_35421_comb + p3_sign_ext_35423_comb;
  assign p3_add_36053_comb = p3_add_35879_comb[31:8] + p2_add_35090[29:6];
  assign p3_add_36055_comb = p3_add_35880_comb[31:8] + p3_sub_35669_comb[31:8];
  assign p3_add_36057_comb = p3_add_35881_comb[31:8] + p3_sub_35672_comb[31:8];
  assign p3_add_36059_comb = p3_add_35882_comb[31:8] + p2_bit_slice_35116;
  assign p3_add_36061_comb = p3_add_35883_comb[31:8] + p2_bit_slice_35119;
  assign p3_add_36063_comb = p3_add_35884_comb[31:8] + p3_sub_35675_comb[31:8];
  assign p3_add_36065_comb = p3_add_35885_comb[31:8] + p3_sub_35678_comb[31:8];
  assign p3_add_36067_comb = p3_add_35886_comb[31:8] + p2_bit_slice_35122;
  assign p3_add_36069_comb = {p3_add_35887_comb, p3_sub_35646_comb[15:11]} + p2_add_35061[29:6];
  assign p3_add_36070_comb = p3_sign_ext_35889_comb[31:8] + p2_add_35090[29:6];
  assign p3_add_36072_comb = {p3_add_35890_comb, p3_sub_35647_comb[15:11]} + p3_sub_35630_comb[31:8];
  assign p3_add_36073_comb = p3_sign_ext_35892_comb[31:8] + p3_sub_35669_comb[31:8];
  assign p3_add_36075_comb = {p3_add_35893_comb, p3_sub_35649_comb[15:11]} + p3_sub_35633_comb[31:8];
  assign p3_add_36076_comb = p3_sign_ext_35895_comb[31:8] + p3_sub_35672_comb[31:8];
  assign p3_add_36078_comb = {p3_add_35896_comb, p2_sub_35078[15:11]} + p2_bit_slice_35154;
  assign p3_add_36079_comb = p3_sign_ext_35898_comb[31:8] + p2_bit_slice_35116;
  assign p3_add_36081_comb = {p3_add_35899_comb, p2_sub_35080[15:11]} + p2_bit_slice_35155;
  assign p3_add_36082_comb = p3_sign_ext_35901_comb[31:8] + p2_bit_slice_35119;
  assign p3_add_36084_comb = {p3_add_35902_comb, p3_sub_35651_comb[15:11]} + p3_sub_35636_comb[31:8];
  assign p3_add_36085_comb = p3_sign_ext_35904_comb[31:8] + p3_sub_35675_comb[31:8];
  assign p3_add_36087_comb = {p3_add_35905_comb, p3_sub_35653_comb[15:11]} + p3_sub_35639_comb[31:8];
  assign p3_add_36088_comb = p3_sign_ext_35907_comb[31:8] + p3_sub_35678_comb[31:8];
  assign p3_add_36090_comb = {p3_add_35908_comb, p2_sub_35082[15:11]} + p2_bit_slice_35156;
  assign p3_add_36091_comb = p3_sign_ext_35910_comb[31:8] + p2_bit_slice_35122;
  assign p3_concat_36093_comb = {p3_add_35984_comb, p3_add_35703_comb[5:0], p3_add_35543_comb[2:1]};
  assign p3_add_36094_comb = p3_sign_ext_35410_comb + p3_sign_ext_35408_comb;
  assign p3_concat_36095_comb = {p3_add_35986_comb, p3_add_35705_comb[5:0], p3_add_35546_comb[2:1]};
  assign p3_add_36096_comb = p3_sign_ext_35414_comb + p3_sign_ext_35412_comb;
  assign p3_concat_36097_comb = {p3_add_35988_comb, p3_add_35707_comb[5:0], p3_add_35551_comb[2:1]};
  assign p3_add_36098_comb = p3_sign_ext_35418_comb + p3_sign_ext_35416_comb;
  assign p3_concat_36099_comb = {p3_add_35990_comb, p3_add_35709_comb[5:0], p3_add_35556_comb[2:1]};
  assign p3_add_36100_comb = p3_sign_ext_35422_comb + p3_sign_ext_35420_comb;
  assign p3_concat_36101_comb = {p3_add_35992_comb, p3_add_35711_comb[5:0], p3_add_35561_comb[2:1]};
  assign p3_sub_36126_comb = {p3_add_35912_comb, 8'h00} - p3_sign_ext_35835_comb;
  assign p3_sub_36127_comb = {p3_add_35914_comb, 8'h00} - p3_sign_ext_35837_comb;
  assign p3_sub_36128_comb = {p3_add_35916_comb, 8'h00} - p3_sign_ext_35839_comb;
  assign p3_sub_36129_comb = {p3_add_35918_comb, 8'h00} - p3_sign_ext_35841_comb;
  assign p3_sub_36130_comb = {p3_add_35920_comb, 8'h00} - p3_sign_ext_35843_comb;
  assign p3_add_36132_comb = p3_sign_ext_35835_comb + p2_add_35172;
  assign p3_add_36134_comb = p3_sign_ext_35837_comb + p3_add_36043_comb;
  assign p3_add_36136_comb = p3_sign_ext_35839_comb + p3_add_36046_comb;
  assign p3_add_36138_comb = p3_sign_ext_35841_comb + p3_add_36049_comb;
  assign p3_add_36140_comb = p3_sign_ext_35843_comb + p3_add_36052_comb;
  assign p3_add_36165_comb = p2_add_35182 + p3_concat_36093_comb;
  assign p3_add_36166_comb = p3_add_36094_comb + p3_concat_36095_comb;
  assign p3_add_36167_comb = p3_add_36096_comb + p3_concat_36097_comb;
  assign p3_add_36168_comb = p3_add_36098_comb + p3_concat_36099_comb;
  assign p3_add_36169_comb = p3_add_36100_comb + p3_concat_36101_comb;
  assign p3_add_36170_comb = p3_sign_ext_35889_comb + {p3_add_35994_comb, p3_sub_35646_comb[10:3]};
  assign p3_add_36171_comb = p3_sign_ext_35892_comb + {p3_add_35996_comb, p3_sub_35647_comb[10:3]};
  assign p3_add_36172_comb = p3_sign_ext_35895_comb + {p3_add_35998_comb, p3_sub_35649_comb[10:3]};
  assign p3_add_36173_comb = p3_sign_ext_35898_comb + {p3_add_36000_comb, p2_sub_35078[10:3]};
  assign p3_add_36174_comb = p3_sign_ext_35901_comb + {p3_add_36002_comb, p2_sub_35080[10:3]};
  assign p3_add_36175_comb = p3_sign_ext_35904_comb + {p3_add_36004_comb, p3_sub_35651_comb[10:3]};
  assign p3_add_36176_comb = p3_sign_ext_35907_comb + {p3_add_36006_comb, p3_sub_35653_comb[10:3]};
  assign p3_add_36177_comb = p3_sign_ext_35910_comb + {p3_add_36008_comb, p2_sub_35082[10:3]};
  assign p3_sub_36178_comb = {p3_add_36010_comb, p2_add_35073[8:1]} - {p3_add_36012_comb, p3_sub_35646_comb[10:3]};
  assign p3_sub_36179_comb = {p3_add_36013_comb, p3_add_35642_comb[8:1]} - {p3_add_36015_comb, p3_sub_35647_comb[10:3]};
  assign p3_sub_36180_comb = {p3_add_36016_comb, p3_add_35643_comb[8:1]} - {p3_add_36018_comb, p3_sub_35649_comb[10:3]};
  assign p3_sub_36181_comb = {p3_add_36019_comb, p2_add_35074[8:1]} - {p3_add_36021_comb, p2_sub_35078[10:3]};
  assign p3_sub_36182_comb = {p3_add_36022_comb, p2_add_35075[8:1]} - {p3_add_36024_comb, p2_sub_35080[10:3]};
  assign p3_sub_36183_comb = {p3_add_36025_comb, p3_add_35644_comb[8:1]} - {p3_add_36027_comb, p3_sub_35651_comb[10:3]};
  assign p3_sub_36184_comb = {p3_add_36028_comb, p3_add_35645_comb[8:1]} - {p3_add_36030_comb, p3_sub_35653_comb[10:3]};
  assign p3_sub_36185_comb = {p3_add_36031_comb, p2_add_35076[8:1]} - {p3_add_36033_comb, p2_sub_35082[10:3]};
  assign p3_add_36186_comb = p3_sub_36126_comb + p2_add_35172;
  assign p3_add_36187_comb = p3_sub_36127_comb + p3_add_36043_comb;
  assign p3_add_36188_comb = p3_sub_36128_comb + p3_add_36046_comb;
  assign p3_add_36189_comb = p3_sub_36129_comb + p3_add_36049_comb;
  assign p3_add_36190_comb = p3_sub_36130_comb + p3_add_36052_comb;
  assign p3_sub_36191_comb = {p3_add_36039_comb, 8'h00} - p3_add_36132_comb;
  assign p3_sub_36192_comb = {p3_add_36041_comb, 8'h00} - p3_add_36134_comb;
  assign p3_sub_36193_comb = {p3_add_36044_comb, 8'h00} - p3_add_36136_comb;
  assign p3_sub_36194_comb = {p3_add_36047_comb, 8'h00} - p3_add_36138_comb;
  assign p3_sub_36195_comb = {p3_add_36050_comb, 8'h00} - p3_add_36140_comb;
  assign p3_sub_36196_comb = p3_concat_35769_comb - {p3_add_36053_comb, p3_add_35879_comb[7:0]};
  assign p3_sub_36197_comb = p3_concat_35771_comb - {p3_add_36055_comb, p3_add_35880_comb[7:0]};
  assign p3_sub_36198_comb = p3_concat_35773_comb - {p3_add_36057_comb, p3_add_35881_comb[7:0]};
  assign p3_sub_36199_comb = p3_concat_35775_comb - {p3_add_36059_comb, p3_add_35882_comb[7:0]};
  assign p3_sub_36200_comb = p3_concat_35777_comb - {p3_add_36061_comb, p3_add_35883_comb[7:0]};
  assign p3_sub_36201_comb = p3_concat_35779_comb - {p3_add_36063_comb, p3_add_35884_comb[7:0]};
  assign p3_sub_36202_comb = p3_concat_35781_comb - {p3_add_36065_comb, p3_add_35885_comb[7:0]};
  assign p3_sub_36203_comb = p3_concat_35783_comb - {p3_add_36067_comb, p3_add_35886_comb[7:0]};
  assign p3_sub_36204_comb = {p3_add_36069_comb, p3_sub_35646_comb[10:3]} - {p3_add_36070_comb, p2_add_35123[8:1]};
  assign p3_sub_36205_comb = {p3_add_36072_comb, p3_sub_35647_comb[10:3]} - {p3_add_36073_comb, p3_add_35754_comb[8:1]};
  assign p3_sub_36206_comb = {p3_add_36075_comb, p3_sub_35649_comb[10:3]} - {p3_add_36076_comb, p3_add_35756_comb[8:1]};
  assign p3_sub_36207_comb = {p3_add_36078_comb, p2_sub_35078[10:3]} - {p3_add_36079_comb, p2_add_35124[8:1]};
  assign p3_sub_36208_comb = {p3_add_36081_comb, p2_sub_35080[10:3]} - {p3_add_36082_comb, p2_add_35125[8:1]};
  assign p3_sub_36209_comb = {p3_add_36084_comb, p3_sub_35651_comb[10:3]} - {p3_add_36085_comb, p3_add_35760_comb[8:1]};
  assign p3_sub_36210_comb = {p3_add_36087_comb, p3_sub_35653_comb[10:3]} - {p3_add_36088_comb, p3_add_35762_comb[8:1]};
  assign p3_sub_36211_comb = {p3_add_36090_comb, p2_sub_35082[10:3]} - {p3_add_36091_comb, p2_add_35126[8:1]};
  assign p3_sub_36212_comb = p3_concat_36093_comb - p2_add_35182;
  assign p3_sub_36213_comb = p3_concat_36095_comb - p3_add_36094_comb;
  assign p3_sub_36214_comb = p3_concat_36097_comb - p3_add_36096_comb;
  assign p3_sub_36215_comb = p3_concat_36099_comb - p3_add_36098_comb;
  assign p3_sub_36216_comb = p3_concat_36101_comb - p3_add_36100_comb;
  assign p3_bit_slice_36217_comb = p3_add_36165_comb[31:14];
  assign p3_bit_slice_36218_comb = p3_add_36166_comb[31:14];
  assign p3_bit_slice_36219_comb = p3_add_36167_comb[31:14];
  assign p3_bit_slice_36220_comb = p3_add_36168_comb[31:14];
  assign p3_bit_slice_36221_comb = p3_add_36169_comb[31:14];
  assign p3_bit_slice_36222_comb = p3_add_36170_comb[31:14];
  assign p3_bit_slice_36223_comb = p3_add_36171_comb[31:14];
  assign p3_bit_slice_36224_comb = p3_add_36172_comb[31:14];
  assign p3_bit_slice_36225_comb = p3_add_36173_comb[31:14];
  assign p3_bit_slice_36226_comb = p3_add_36174_comb[31:14];
  assign p3_bit_slice_36227_comb = p3_add_36175_comb[31:14];
  assign p3_bit_slice_36228_comb = p3_add_36176_comb[31:14];
  assign p3_bit_slice_36229_comb = p3_add_36177_comb[31:14];
  assign p3_bit_slice_36230_comb = p3_sub_36178_comb[31:14];
  assign p3_bit_slice_36231_comb = p3_sub_36179_comb[31:14];
  assign p3_bit_slice_36232_comb = p3_sub_36180_comb[31:14];
  assign p3_bit_slice_36233_comb = p3_sub_36181_comb[31:14];
  assign p3_bit_slice_36234_comb = p3_sub_36182_comb[31:14];
  assign p3_bit_slice_36235_comb = p3_sub_36183_comb[31:14];
  assign p3_bit_slice_36236_comb = p3_sub_36184_comb[31:14];
  assign p3_bit_slice_36237_comb = p3_sub_36185_comb[31:14];
  assign p3_bit_slice_36238_comb = p3_add_36186_comb[31:14];
  assign p3_bit_slice_36239_comb = p3_add_36187_comb[31:14];
  assign p3_bit_slice_36240_comb = p3_add_36188_comb[31:14];
  assign p3_bit_slice_36241_comb = p3_add_36189_comb[31:14];
  assign p3_bit_slice_36242_comb = p3_add_36190_comb[31:14];
  assign p3_bit_slice_36243_comb = p3_sub_36191_comb[31:14];
  assign p3_bit_slice_36244_comb = p3_sub_36192_comb[31:14];
  assign p3_bit_slice_36245_comb = p3_sub_36193_comb[31:14];
  assign p3_bit_slice_36246_comb = p3_sub_36194_comb[31:14];
  assign p3_bit_slice_36247_comb = p3_sub_36195_comb[31:14];
  assign p3_bit_slice_36248_comb = p3_sub_36196_comb[31:14];
  assign p3_bit_slice_36249_comb = p3_sub_36197_comb[31:14];
  assign p3_bit_slice_36250_comb = p3_sub_36198_comb[31:14];
  assign p3_bit_slice_36251_comb = p3_sub_36199_comb[31:14];
  assign p3_bit_slice_36252_comb = p3_sub_36200_comb[31:14];
  assign p3_bit_slice_36253_comb = p3_sub_36201_comb[31:14];
  assign p3_bit_slice_36254_comb = p3_sub_36202_comb[31:14];
  assign p3_bit_slice_36255_comb = p3_sub_36203_comb[31:14];
  assign p3_bit_slice_36256_comb = p3_sub_36204_comb[31:14];
  assign p3_bit_slice_36257_comb = p3_sub_36205_comb[31:14];
  assign p3_bit_slice_36258_comb = p3_sub_36206_comb[31:14];
  assign p3_bit_slice_36259_comb = p3_sub_36207_comb[31:14];
  assign p3_bit_slice_36260_comb = p3_sub_36208_comb[31:14];
  assign p3_bit_slice_36261_comb = p3_sub_36209_comb[31:14];
  assign p3_bit_slice_36262_comb = p3_sub_36210_comb[31:14];
  assign p3_bit_slice_36263_comb = p3_sub_36211_comb[31:14];
  assign p3_bit_slice_36264_comb = p3_sub_36212_comb[31:14];
  assign p3_bit_slice_36265_comb = p3_sub_36213_comb[31:14];
  assign p3_bit_slice_36266_comb = p3_sub_36214_comb[31:14];
  assign p3_bit_slice_36267_comb = p3_sub_36215_comb[31:14];
  assign p3_bit_slice_36268_comb = p3_sub_36216_comb[31:14];
  assign p3_array_36333_comb[0] = {{14{p3_bit_slice_36217_comb[17]}}, p3_bit_slice_36217_comb};
  assign p3_array_36333_comb[1] = {{14{p3_bit_slice_36218_comb[17]}}, p3_bit_slice_36218_comb};
  assign p3_array_36333_comb[2] = {{14{p3_bit_slice_36219_comb[17]}}, p3_bit_slice_36219_comb};
  assign p3_array_36333_comb[3] = {{14{p2_bit_slice_35210[17]}}, p2_bit_slice_35210};
  assign p3_array_36333_comb[4] = {{14{p2_bit_slice_35211[17]}}, p2_bit_slice_35211};
  assign p3_array_36333_comb[5] = {{14{p3_bit_slice_36220_comb[17]}}, p3_bit_slice_36220_comb};
  assign p3_array_36333_comb[6] = {{14{p3_bit_slice_36221_comb[17]}}, p3_bit_slice_36221_comb};
  assign p3_array_36333_comb[7] = {{14{p2_bit_slice_35212[17]}}, p2_bit_slice_35212};
  assign p3_array_36333_comb[8] = {{14{p3_bit_slice_36222_comb[17]}}, p3_bit_slice_36222_comb};
  assign p3_array_36333_comb[9] = {{14{p3_bit_slice_36223_comb[17]}}, p3_bit_slice_36223_comb};
  assign p3_array_36333_comb[10] = {{14{p3_bit_slice_36224_comb[17]}}, p3_bit_slice_36224_comb};
  assign p3_array_36333_comb[11] = {{14{p3_bit_slice_36225_comb[17]}}, p3_bit_slice_36225_comb};
  assign p3_array_36333_comb[12] = {{14{p3_bit_slice_36226_comb[17]}}, p3_bit_slice_36226_comb};
  assign p3_array_36333_comb[13] = {{14{p3_bit_slice_36227_comb[17]}}, p3_bit_slice_36227_comb};
  assign p3_array_36333_comb[14] = {{14{p3_bit_slice_36228_comb[17]}}, p3_bit_slice_36228_comb};
  assign p3_array_36333_comb[15] = {{14{p3_bit_slice_36229_comb[17]}}, p3_bit_slice_36229_comb};
  assign p3_array_36333_comb[16] = {{14{p3_bit_slice_36230_comb[17]}}, p3_bit_slice_36230_comb};
  assign p3_array_36333_comb[17] = {{14{p3_bit_slice_36231_comb[17]}}, p3_bit_slice_36231_comb};
  assign p3_array_36333_comb[18] = {{14{p3_bit_slice_36232_comb[17]}}, p3_bit_slice_36232_comb};
  assign p3_array_36333_comb[19] = {{14{p3_bit_slice_36233_comb[17]}}, p3_bit_slice_36233_comb};
  assign p3_array_36333_comb[20] = {{14{p3_bit_slice_36234_comb[17]}}, p3_bit_slice_36234_comb};
  assign p3_array_36333_comb[21] = {{14{p3_bit_slice_36235_comb[17]}}, p3_bit_slice_36235_comb};
  assign p3_array_36333_comb[22] = {{14{p3_bit_slice_36236_comb[17]}}, p3_bit_slice_36236_comb};
  assign p3_array_36333_comb[23] = {{14{p3_bit_slice_36237_comb[17]}}, p3_bit_slice_36237_comb};
  assign p3_array_36333_comb[24] = {{14{p3_bit_slice_36238_comb[17]}}, p3_bit_slice_36238_comb};
  assign p3_array_36333_comb[25] = {{14{p3_bit_slice_36239_comb[17]}}, p3_bit_slice_36239_comb};
  assign p3_array_36333_comb[26] = {{14{p3_bit_slice_36240_comb[17]}}, p3_bit_slice_36240_comb};
  assign p3_array_36333_comb[27] = {{14{p2_bit_slice_35213[17]}}, p2_bit_slice_35213};
  assign p3_array_36333_comb[28] = {{14{p2_bit_slice_35214[17]}}, p2_bit_slice_35214};
  assign p3_array_36333_comb[29] = {{14{p3_bit_slice_36241_comb[17]}}, p3_bit_slice_36241_comb};
  assign p3_array_36333_comb[30] = {{14{p3_bit_slice_36242_comb[17]}}, p3_bit_slice_36242_comb};
  assign p3_array_36333_comb[31] = {{14{p2_bit_slice_35215[17]}}, p2_bit_slice_35215};
  assign p3_array_36333_comb[32] = {{14{p3_bit_slice_36243_comb[17]}}, p3_bit_slice_36243_comb};
  assign p3_array_36333_comb[33] = {{14{p3_bit_slice_36244_comb[17]}}, p3_bit_slice_36244_comb};
  assign p3_array_36333_comb[34] = {{14{p3_bit_slice_36245_comb[17]}}, p3_bit_slice_36245_comb};
  assign p3_array_36333_comb[35] = {{14{p2_bit_slice_35216[17]}}, p2_bit_slice_35216};
  assign p3_array_36333_comb[36] = {{14{p2_bit_slice_35217[17]}}, p2_bit_slice_35217};
  assign p3_array_36333_comb[37] = {{14{p3_bit_slice_36246_comb[17]}}, p3_bit_slice_36246_comb};
  assign p3_array_36333_comb[38] = {{14{p3_bit_slice_36247_comb[17]}}, p3_bit_slice_36247_comb};
  assign p3_array_36333_comb[39] = {{14{p2_bit_slice_35218[17]}}, p2_bit_slice_35218};
  assign p3_array_36333_comb[40] = {{14{p3_bit_slice_36248_comb[17]}}, p3_bit_slice_36248_comb};
  assign p3_array_36333_comb[41] = {{14{p3_bit_slice_36249_comb[17]}}, p3_bit_slice_36249_comb};
  assign p3_array_36333_comb[42] = {{14{p3_bit_slice_36250_comb[17]}}, p3_bit_slice_36250_comb};
  assign p3_array_36333_comb[43] = {{14{p3_bit_slice_36251_comb[17]}}, p3_bit_slice_36251_comb};
  assign p3_array_36333_comb[44] = {{14{p3_bit_slice_36252_comb[17]}}, p3_bit_slice_36252_comb};
  assign p3_array_36333_comb[45] = {{14{p3_bit_slice_36253_comb[17]}}, p3_bit_slice_36253_comb};
  assign p3_array_36333_comb[46] = {{14{p3_bit_slice_36254_comb[17]}}, p3_bit_slice_36254_comb};
  assign p3_array_36333_comb[47] = {{14{p3_bit_slice_36255_comb[17]}}, p3_bit_slice_36255_comb};
  assign p3_array_36333_comb[48] = {{14{p3_bit_slice_36256_comb[17]}}, p3_bit_slice_36256_comb};
  assign p3_array_36333_comb[49] = {{14{p3_bit_slice_36257_comb[17]}}, p3_bit_slice_36257_comb};
  assign p3_array_36333_comb[50] = {{14{p3_bit_slice_36258_comb[17]}}, p3_bit_slice_36258_comb};
  assign p3_array_36333_comb[51] = {{14{p3_bit_slice_36259_comb[17]}}, p3_bit_slice_36259_comb};
  assign p3_array_36333_comb[52] = {{14{p3_bit_slice_36260_comb[17]}}, p3_bit_slice_36260_comb};
  assign p3_array_36333_comb[53] = {{14{p3_bit_slice_36261_comb[17]}}, p3_bit_slice_36261_comb};
  assign p3_array_36333_comb[54] = {{14{p3_bit_slice_36262_comb[17]}}, p3_bit_slice_36262_comb};
  assign p3_array_36333_comb[55] = {{14{p3_bit_slice_36263_comb[17]}}, p3_bit_slice_36263_comb};
  assign p3_array_36333_comb[56] = {{14{p3_bit_slice_36264_comb[17]}}, p3_bit_slice_36264_comb};
  assign p3_array_36333_comb[57] = {{14{p3_bit_slice_36265_comb[17]}}, p3_bit_slice_36265_comb};
  assign p3_array_36333_comb[58] = {{14{p3_bit_slice_36266_comb[17]}}, p3_bit_slice_36266_comb};
  assign p3_array_36333_comb[59] = {{14{p2_bit_slice_35219[17]}}, p2_bit_slice_35219};
  assign p3_array_36333_comb[60] = {{14{p2_bit_slice_35220[17]}}, p2_bit_slice_35220};
  assign p3_array_36333_comb[61] = {{14{p3_bit_slice_36267_comb[17]}}, p3_bit_slice_36267_comb};
  assign p3_array_36333_comb[62] = {{14{p3_bit_slice_36268_comb[17]}}, p3_bit_slice_36268_comb};
  assign p3_array_36333_comb[63] = {{14{p2_bit_slice_35221[17]}}, p2_bit_slice_35221};

  // Registers for pipe stage 3:
  reg [31:0] p3_array_36333[64];
  always_ff @ (posedge clk) begin
    p3_array_36333 <= p3_array_36333_comb;
  end
  assign out = {p3_array_36333[63], p3_array_36333[62], p3_array_36333[61], p3_array_36333[60], p3_array_36333[59], p3_array_36333[58], p3_array_36333[57], p3_array_36333[56], p3_array_36333[55], p3_array_36333[54], p3_array_36333[53], p3_array_36333[52], p3_array_36333[51], p3_array_36333[50], p3_array_36333[49], p3_array_36333[48], p3_array_36333[47], p3_array_36333[46], p3_array_36333[45], p3_array_36333[44], p3_array_36333[43], p3_array_36333[42], p3_array_36333[41], p3_array_36333[40], p3_array_36333[39], p3_array_36333[38], p3_array_36333[37], p3_array_36333[36], p3_array_36333[35], p3_array_36333[34], p3_array_36333[33], p3_array_36333[32], p3_array_36333[31], p3_array_36333[30], p3_array_36333[29], p3_array_36333[28], p3_array_36333[27], p3_array_36333[26], p3_array_36333[25], p3_array_36333[24], p3_array_36333[23], p3_array_36333[22], p3_array_36333[21], p3_array_36333[20], p3_array_36333[19], p3_array_36333[18], p3_array_36333[17], p3_array_36333[16], p3_array_36333[15], p3_array_36333[14], p3_array_36333[13], p3_array_36333[12], p3_array_36333[11], p3_array_36333[10], p3_array_36333[9], p3_array_36333[8], p3_array_36333[7], p3_array_36333[6], p3_array_36333[5], p3_array_36333[4], p3_array_36333[3], p3_array_36333[2], p3_array_36333[1], p3_array_36333[0]};
endmodule
